--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- Written by build_rom.py for project 'cpu_test'.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.light52_pkg.all;

package obj_code_pkg is

-- Size of XCODE memory in bytes.
constant XCODE_SIZE : natural := 40000;
-- Size of XDATA memory in bytes.
constant XDATA_SIZE : natural := 512;

-- Object code initialization constant.
constant object_code : t_obj_code(0 to 32800) := (
    X"02", X"00", X"30", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"75", X"6e", X"00", X"75", X"99", X"41", X"75", X"99", 
    X"61", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"99", X"62", X"80", X"05", X"75", X"99", 
    X"63", X"80", X"18", X"75", X"e0", X"5a", X"b4", X"5a", 
    X"f5", X"b4", X"7a", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"b4", X"7a", X"e9", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"75", X"60", X"02", X"d5", X"60", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"d5", 
    X"60", X"05", X"75", X"99", X"64", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"60", X"a5", 
    X"e5", X"60", X"b4", X"a5", X"05", X"75", X"99", X"65", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", X"99", 
    X"42", X"78", X"81", X"e8", X"b4", X"81", X"2f", X"79", 
    X"43", X"e9", X"b4", X"43", X"29", X"7a", X"27", X"ea", 
    X"b4", X"27", X"23", X"7b", X"c2", X"eb", X"b4", X"c2", 
    X"1d", X"7c", X"f1", X"ec", X"b4", X"f1", X"17", X"7d", 
    X"04", X"ed", X"b4", X"04", X"11", X"7e", X"92", X"ee", 
    X"b4", X"92", X"0b", X"7f", X"1f", X"ef", X"b4", X"1f", 
    X"05", X"75", X"99", X"61", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"d0", X"80", X"40", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"50", 
    X"07", X"75", X"d0", X"00", X"40", X"02", X"50", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", 
    X"62", X"78", X"92", X"b8", X"91", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"78", X"91", X"b8", X"91", 
    X"fb", X"79", X"a3", X"b9", X"a2", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"79", X"a2", X"b9", X"a2", 
    X"fb", X"7a", X"b4", X"ba", X"b3", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7a", X"b3", X"ba", X"b3", 
    X"fb", X"7b", X"c5", X"bb", X"c4", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7b", X"c4", X"bb", X"c4", 
    X"fb", X"7c", X"d6", X"bc", X"d5", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7c", X"d5", X"bc", X"d5", 
    X"fb", X"7d", X"e7", X"bd", X"e6", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7d", X"e6", X"bd", X"e6", 
    X"fb", X"7e", X"f8", X"be", X"f7", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7e", X"f7", X"be", X"f7", 
    X"fb", X"7f", X"09", X"bf", X"08", X"08", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7f", X"08", X"bf", X"08", 
    X"fb", X"75", X"d0", X"00", X"78", X"34", X"b8", X"35", 
    X"00", X"50", X"0f", X"b8", X"34", X"00", X"40", X"0a", 
    X"b8", X"33", X"00", X"40", X"05", X"75", X"99", X"63", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"75", X"d0", X"80", X"c3", X"40", X"0b", X"d3", X"50", 
    X"08", X"b3", X"40", X"05", X"75", X"99", X"64", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"78", 
    X"60", X"75", X"60", X"12", X"e5", X"60", X"b4", X"12", 
    X"1d", X"76", X"f5", X"e5", X"60", X"b4", X"f5", X"16", 
    X"79", X"60", X"75", X"60", X"12", X"e5", X"60", X"b4", 
    X"12", X"0c", X"77", X"f5", X"e5", X"60", X"b4", X"f5", 
    X"05", X"75", X"99", X"65", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"78", X"30", X"76", X"13", 
    X"b6", X"12", X"08", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"76", X"12", X"b6", X"12", X"fb", X"79", X"30", 
    X"77", X"35", X"b7", X"34", X"08", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"77", X"34", X"b7", X"34", X"fb", 
    X"78", X"30", X"c3", X"76", X"34", X"b6", X"35", X"00", 
    X"50", X"0f", X"b6", X"34", X"00", X"40", X"0a", X"b6", 
    X"33", X"00", X"40", X"05", X"75", X"99", X"66", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"60", X"c0", X"75", X"31", X"c1", X"75", X"32", X"c2", 
    X"c3", X"74", X"c1", X"b5", X"31", X"1d", X"40", X"1b", 
    X"b5", X"32", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"50", X"10", X"b5", X"60", X"06", X"75", X"99", 
    X"24", X"75", X"6e", X"01", X"40", X"05", X"75", X"99", 
    X"67", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"60", X"c0", X"75", X"f0", X"c1", X"75", 
    X"32", X"c2", X"c3", X"74", X"c1", X"78", X"42", X"b5", 
    X"f0", X"1d", X"40", X"1b", X"b5", X"32", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"50", X"10", X"b5", 
    X"60", X"06", X"75", X"99", X"24", X"75", X"6e", X"01", 
    X"40", X"05", X"75", X"99", X"68", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", X"0d", 
    X"75", X"99", X"0a", X"75", X"99", X"43", X"75", X"2f", 
    X"80", X"80", X"0e", X"30", X"7f", X"1c", X"30", X"7e", 
    X"11", X"75", X"99", X"3f", X"75", X"6e", X"01", X"80", 
    X"11", X"20", X"7f", X"ef", X"75", X"99", X"21", X"75", 
    X"6e", X"01", X"20", X"7e", X"05", X"75", X"99", X"61", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"75", X"e0", X"79", X"b4", X"79", X"0a", X"74", X"5a", 
    X"b4", X"5a", X"05", X"75", X"99", X"62", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"74", X"80", 
    X"80", X"0e", X"60", X"1b", X"74", X"00", X"60", X"10", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"80", X"0f", 
    X"70", X"f0", X"75", X"99", X"21", X"75", X"6e", X"01", 
    X"70", X"05", X"75", X"99", X"63", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"2f", X"80", 
    X"20", X"7f", X"02", X"80", X"0f", X"c2", X"7f", X"20", 
    X"7f", X"0a", X"b2", X"7f", X"30", X"7f", X"05", X"75", 
    X"99", X"64", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"2e", X"08", X"c3", X"82", X"73", 
    X"40", X"1f", X"d3", X"82", X"73", X"50", X"1a", X"b0", 
    X"72", X"50", X"16", X"72", X"73", X"50", X"12", X"72", 
    X"72", X"50", X"0e", X"c3", X"72", X"73", X"50", X"09", 
    X"a0", X"72", X"50", X"05", X"75", X"99", X"65", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"2e", X"08", X"c3", X"a2", X"73", X"50", X"15", X"a2", 
    X"72", X"40", X"11", X"c3", X"92", X"71", X"20", X"71", 
    X"0b", X"d3", X"92", X"71", X"30", X"71", X"05", X"75", 
    X"99", X"66", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"2e", X"00", X"d2", X"73", X"a2", 
    X"73", X"50", X"0b", X"d2", X"72", X"a2", X"72", X"50", 
    X"05", X"75", X"99", X"67", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"2e", X"08", X"80", 
    X"09", X"a2", X"73", X"40", X"0f", X"10", X"72", X"0c", 
    X"80", X"05", X"10", X"73", X"f4", X"80", X"05", X"75", 
    X"99", X"68", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"2f", X"00", X"75", X"f0", X"80", 
    X"80", X"0e", X"30", X"f7", X"1c", X"30", X"f6", X"11", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"80", X"11", 
    X"20", X"f7", X"ef", X"75", X"99", X"21", X"75", X"6e", 
    X"01", X"20", X"f6", X"05", X"75", X"99", X"69", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"f0", X"80", X"20", X"f7", X"02", X"80", X"0f", X"c2", 
    X"f7", X"20", X"f7", X"0a", X"b2", X"f7", X"30", X"f7", 
    X"05", X"75", X"99", X"6a", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"f0", X"08", X"c3", 
    X"82", X"f3", X"40", X"1f", X"d3", X"82", X"f3", X"50", 
    X"1a", X"b0", X"f2", X"50", X"16", X"72", X"f3", X"50", 
    X"12", X"72", X"f2", X"50", X"0e", X"c3", X"72", X"f3", 
    X"50", X"09", X"a0", X"f2", X"50", X"05", X"75", X"99", 
    X"6b", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"f0", X"08", X"c3", X"a2", X"f3", X"50", 
    X"15", X"a2", X"f2", X"40", X"11", X"c3", X"92", X"f1", 
    X"20", X"f1", X"0b", X"d3", X"92", X"f1", X"30", X"f1", 
    X"05", X"75", X"99", X"6c", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"2e", X"00", X"d2", 
    X"f3", X"a2", X"f3", X"50", X"0b", X"d2", X"f2", X"a2", 
    X"f2", X"50", X"05", X"75", X"99", X"6d", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"f0", 
    X"08", X"80", X"09", X"a2", X"f3", X"40", X"0f", X"10", 
    X"f2", X"0c", X"80", X"05", X"10", X"f3", X"f4", X"80", 
    X"05", X"75", X"99", X"6e", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"e0", X"08", X"80", 
    X"09", X"a2", X"e3", X"40", X"0f", X"10", X"e2", X"0c", 
    X"80", X"05", X"10", X"e3", X"f4", X"80", X"05", X"75", 
    X"99", X"6f", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"2e", X"00", X"d2", X"e3", X"a2", 
    X"e3", X"50", X"0b", X"d2", X"e2", X"a2", X"e2", X"50", 
    X"05", X"75", X"99", X"70", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"e0", X"80", X"20", 
    X"e7", X"02", X"80", X"0f", X"c2", X"e7", X"20", X"e7", 
    X"0a", X"b2", X"e7", X"30", X"e7", X"05", X"75", X"99", 
    X"71", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", 
    X"99", X"44", X"74", X"85", X"64", X"44", X"60", X"09", 
    X"64", X"c1", X"70", X"05", X"75", X"99", X"61", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"74", 
    X"85", X"00", X"c3", X"33", X"f5", X"60", X"64", X"0a", 
    X"70", X"16", X"e5", X"60", X"33", X"64", X"15", X"70", 
    X"0f", X"74", X"85", X"00", X"c3", X"33", X"50", X"08", 
    X"33", X"40", X"05", X"75", X"99", X"62", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"74", X"85", 
    X"c3", X"13", X"f5", X"60", X"00", X"64", X"42", X"70", 
    X"15", X"e5", X"60", X"13", X"64", X"a1", X"70", X"0e", 
    X"74", X"85", X"c3", X"13", X"50", X"08", X"13", X"40", 
    X"05", X"75", X"99", X"63", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"74", X"85", X"c3", X"23", 
    X"f5", X"60", X"64", X"0b", X"70", X"28", X"e5", X"60", 
    X"d3", X"23", X"64", X"16", X"70", X"20", X"74", X"85", 
    X"c3", X"03", X"f5", X"60", X"64", X"c2", X"70", X"16", 
    X"e5", X"60", X"03", X"64", X"61", X"70", X"0f", X"74", 
    X"ff", X"c3", X"23", X"40", X"09", X"03", X"03", X"40", 
    X"05", X"75", X"99", X"64", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"99", X"0d", X"75", 
    X"99", X"0a", X"75", X"99", X"45", X"74", X"80", X"04", 
    X"b4", X"81", X"0e", X"74", X"ff", X"c3", X"04", X"40", 
    X"08", X"b4", X"00", X"05", X"75", X"99", X"61", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"78", 
    X"66", X"78", X"80", X"08", X"b8", X"81", X"77", X"78", 
    X"ff", X"c3", X"08", X"40", X"71", X"b8", X"00", X"6e", 
    X"79", X"80", X"09", X"b9", X"81", X"68", X"79", X"ff", 
    X"c3", X"09", X"40", X"62", X"b9", X"00", X"5f", X"7a", 
    X"80", X"0a", X"ba", X"81", X"59", X"7a", X"ff", X"c3", 
    X"0a", X"40", X"53", X"ba", X"00", X"50", X"7b", X"80", 
    X"0b", X"bb", X"81", X"4a", X"7b", X"ff", X"c3", X"0b", 
    X"40", X"44", X"bb", X"00", X"41", X"7c", X"80", X"0c", 
    X"bc", X"81", X"3b", X"7c", X"ff", X"c3", X"0c", X"40", 
    X"35", X"bc", X"00", X"32", X"7d", X"80", X"0d", X"bd", 
    X"81", X"2c", X"7d", X"ff", X"c3", X"0d", X"40", X"26", 
    X"bd", X"00", X"23", X"7e", X"80", X"0e", X"be", X"81", 
    X"1d", X"7e", X"ff", X"c3", X"0e", X"40", X"17", X"be", 
    X"00", X"14", X"7f", X"80", X"0f", X"bf", X"81", X"0e", 
    X"7f", X"ff", X"c3", X"0f", X"40", X"08", X"bf", X"00", 
    X"05", X"75", X"99", X"62", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"78", X"60", X"79", X"31", 
    X"76", X"80", X"06", X"b6", X"81", X"1d", X"76", X"ff", 
    X"c3", X"06", X"40", X"17", X"b6", X"00", X"14", X"77", 
    X"80", X"07", X"b7", X"81", X"0e", X"77", X"ff", X"c3", 
    X"07", X"40", X"08", X"b7", X"00", X"05", X"75", X"99", 
    X"63", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"60", X"34", X"e5", X"60", X"b4", X"34", 
    X"05", X"75", X"99", X"64", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"39", X"80", X"05", 
    X"39", X"e5", X"39", X"b4", X"81", X"29", X"75", X"39", 
    X"ff", X"c3", X"05", X"39", X"40", X"21", X"e5", X"39", 
    X"b4", X"00", X"1c", X"75", X"f0", X"80", X"05", X"f0", 
    X"e5", X"f0", X"b4", X"81", X"12", X"75", X"f0", X"ff", 
    X"c3", X"05", X"f0", X"40", X"0a", X"e5", X"f0", X"b4", 
    X"00", X"05", X"75", X"99", X"65", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"74", X"01", X"14", 
    X"b4", X"00", X"0c", X"c3", X"14", X"40", X"08", X"b4", 
    X"ff", X"05", X"75", X"99", X"66", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"78", X"66", X"78", 
    X"01", X"18", X"b8", X"00", X"67", X"c3", X"18", X"40", 
    X"63", X"b8", X"ff", X"60", X"79", X"01", X"19", X"b9", 
    X"00", X"5a", X"c3", X"19", X"40", X"56", X"b9", X"ff", 
    X"53", X"7a", X"01", X"1a", X"ba", X"00", X"4d", X"c3", 
    X"1a", X"40", X"49", X"ba", X"ff", X"46", X"7b", X"01", 
    X"1b", X"bb", X"00", X"40", X"c3", X"1b", X"40", X"3c", 
    X"bb", X"ff", X"39", X"7c", X"01", X"1c", X"bc", X"00", 
    X"33", X"c3", X"1c", X"40", X"2f", X"bc", X"ff", X"2c", 
    X"7d", X"01", X"1d", X"bd", X"00", X"26", X"c3", X"1d", 
    X"40", X"22", X"bd", X"ff", X"1f", X"7e", X"01", X"1e", 
    X"be", X"00", X"19", X"c3", X"1e", X"40", X"15", X"be", 
    X"ff", X"12", X"7f", X"01", X"1f", X"bf", X"00", X"0c", 
    X"c3", X"1f", X"40", X"08", X"bf", X"ff", X"05", X"75", 
    X"99", X"67", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"78", X"60", X"79", X"31", X"76", X"01", 
    X"16", X"b6", X"00", X"19", X"c3", X"16", X"40", X"15", 
    X"b6", X"ff", X"12", X"77", X"01", X"17", X"b7", X"00", 
    X"0c", X"c3", X"17", X"40", X"08", X"b7", X"ff", X"05", 
    X"75", X"99", X"68", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"75", X"39", X"01", X"15", X"39", 
    X"e5", X"39", X"b4", X"00", X"29", X"75", X"39", X"00", 
    X"c3", X"15", X"39", X"40", X"21", X"e5", X"39", X"b4", 
    X"ff", X"1c", X"75", X"f0", X"01", X"15", X"f0", X"e5", 
    X"f0", X"b4", X"00", X"12", X"75", X"f0", X"00", X"c3", 
    X"15", X"f0", X"40", X"0a", X"e5", X"f0", X"b4", X"ff", 
    X"05", X"75", X"99", X"69", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"99", X"0d", X"75", 
    X"99", X"0a", X"75", X"99", X"46", X"78", X"91", X"88", 
    X"39", X"e5", X"39", X"b4", X"91", X"44", X"79", X"92", 
    X"89", X"39", X"e5", X"39", X"b4", X"92", X"3b", X"7a", 
    X"93", X"8a", X"39", X"e5", X"39", X"b4", X"93", X"32", 
    X"7b", X"94", X"8b", X"39", X"e5", X"39", X"b4", X"94", 
    X"29", X"7c", X"95", X"8c", X"39", X"e5", X"39", X"b4", 
    X"95", X"20", X"7d", X"96", X"8d", X"39", X"e5", X"39", 
    X"b4", X"96", X"17", X"7e", X"97", X"8e", X"39", X"e5", 
    X"39", X"b4", X"97", X"0e", X"7f", X"98", X"8f", X"39", 
    X"e5", X"39", X"b4", X"98", X"05", X"75", X"99", X"61", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"76", X"91", X"86", X"39", X"e5", X"39", X"b4", X"91", 
    X"0e", X"77", X"92", X"87", X"39", X"e5", X"39", X"b4", 
    X"92", X"05", X"75", X"99", X"62", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"31", X"91", 
    X"85", X"31", X"39", X"e5", X"39", X"b4", X"91", X"1b", 
    X"75", X"31", X"91", X"85", X"31", X"f0", X"e5", X"f0", 
    X"b4", X"91", X"10", X"75", X"f0", X"91", X"85", X"f0", 
    X"31", X"e5", X"31", X"b4", X"91", X"05", X"75", X"99", 
    X"63", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"39", X"91", X"a8", X"39", X"b8", X"91", 
    X"3d", X"75", X"39", X"92", X"a9", X"39", X"b9", X"92", 
    X"35", X"75", X"39", X"93", X"aa", X"39", X"ba", X"93", 
    X"2d", X"75", X"39", X"94", X"ab", X"39", X"bb", X"94", 
    X"25", X"75", X"39", X"95", X"ac", X"39", X"bc", X"95", 
    X"1d", X"75", X"39", X"96", X"ad", X"39", X"bd", X"96", 
    X"15", X"75", X"39", X"97", X"ae", X"39", X"be", X"97", 
    X"0d", X"75", X"39", X"98", X"af", X"39", X"bf", X"98", 
    X"05", X"75", X"99", X"64", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"78", X"60", X"79", X"31", 
    X"75", X"39", X"91", X"a6", X"39", X"b6", X"91", X"0d", 
    X"75", X"39", X"92", X"a7", X"39", X"b7", X"92", X"05", 
    X"75", X"99", X"65", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"74", X"91", X"f8", X"b8", X"91", 
    X"2f", X"74", X"92", X"f9", X"b9", X"92", X"29", X"74", 
    X"93", X"fa", X"ba", X"93", X"23", X"74", X"94", X"fb", 
    X"bb", X"94", X"1d", X"74", X"95", X"fc", X"bc", X"95", 
    X"17", X"74", X"96", X"fd", X"bd", X"96", X"11", X"74", 
    X"97", X"fe", X"be", X"97", X"0b", X"74", X"98", X"ff", 
    X"bf", X"98", X"05", X"75", X"99", X"66", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"78", X"60", 
    X"79", X"31", X"74", X"91", X"f6", X"b6", X"91", X"0b", 
    X"74", X"92", X"f7", X"b7", X"92", X"05", X"75", X"99", 
    X"67", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"60", X"79", X"78", X"00", X"74", X"34", 
    X"f5", X"60", X"a8", X"60", X"b8", X"34", X"05", X"75", 
    X"99", X"68", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"74", X"00", X"79", X"31", X"75", X"31", 
    X"56", X"78", X"60", X"75", X"60", X"34", X"e6", X"b4", 
    X"34", X"09", X"e7", X"b4", X"56", X"05", X"75", X"99", 
    X"69", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", 
    X"99", X"47", X"74", X"55", X"e4", X"70", X"11", X"74", 
    X"55", X"f4", X"b4", X"aa", X"0b", X"74", X"97", X"c4", 
    X"b4", X"79", X"05", X"75", X"99", X"61", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"83", 
    X"12", X"75", X"82", X"fd", X"a3", X"e5", X"83", X"b4", 
    X"12", X"20", X"e5", X"82", X"b4", X"fe", X"1b", X"a3", 
    X"e5", X"83", X"b4", X"12", X"15", X"e5", X"82", X"b4", 
    X"ff", X"10", X"a3", X"e5", X"83", X"b4", X"13", X"0a", 
    X"e5", X"82", X"b4", X"00", X"05", X"75", X"99", X"62", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"74", X"34", X"75", X"13", X"57", X"c5", X"13", X"b4", 
    X"57", X"19", X"e5", X"13", X"b4", X"34", X"14", X"74", 
    X"34", X"75", X"f0", X"57", X"c5", X"f0", X"b4", X"57", 
    X"0a", X"e5", X"f0", X"b4", X"34", X"05", X"75", X"99", 
    X"63", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"74", X"91", X"75", X"29", X"78", X"78", X"29", 
    X"c6", X"b4", X"78", X"1a", X"e5", X"29", X"b4", X"91", 
    X"15", X"74", X"92", X"75", X"2a", X"78", X"79", X"2a", 
    X"c7", X"b4", X"78", X"0a", X"e5", X"2a", X"b4", X"92", 
    X"05", X"75", X"99", X"64", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"74", X"d4", X"78", X"55", 
    X"c8", X"b8", X"d4", X"55", X"b4", X"55", X"52", X"74", 
    X"d3", X"79", X"54", X"c9", X"b9", X"d3", X"4a", X"b4", 
    X"54", X"47", X"74", X"d2", X"7a", X"53", X"ca", X"ba", 
    X"d2", X"3f", X"b4", X"53", X"3c", X"74", X"d1", X"7b", 
    X"52", X"cb", X"bb", X"d1", X"34", X"b4", X"52", X"31", 
    X"74", X"d0", X"7c", X"51", X"cc", X"bc", X"d0", X"29", 
    X"b4", X"51", X"26", X"74", X"cf", X"7d", X"50", X"cd", 
    X"bd", X"cf", X"1e", X"b4", X"50", X"1b", X"74", X"ce", 
    X"7e", X"4f", X"ce", X"be", X"ce", X"13", X"b4", X"4f", 
    X"10", X"74", X"cd", X"7f", X"4e", X"cf", X"bf", X"cd", 
    X"08", X"b4", X"4e", X"05", X"75", X"99", X"65", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"99", X"0d", X"75", X"99", X"0a", X"75", X"99", X"48", 
    X"75", X"60", X"3c", X"74", X"99", X"55", X"60", X"b4", 
    X"18", X"29", X"78", X"60", X"76", X"3c", X"74", X"99", 
    X"56", X"b4", X"18", X"1f", X"79", X"31", X"77", X"3c", 
    X"74", X"99", X"57", X"b4", X"18", X"15", X"78", X"3c", 
    X"74", X"99", X"58", X"b4", X"18", X"0d", X"79", X"3c", 
    X"74", X"99", X"59", X"b4", X"18", X"05", X"75", X"99", 
    X"61", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"7a", X"3c", X"74", X"99", X"5a", X"b4", X"18", 
    X"0d", X"7b", X"3c", X"74", X"99", X"5b", X"b4", X"18", 
    X"05", X"75", X"99", X"62", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7c", X"3c", X"74", X"99", 
    X"5c", X"b4", X"18", X"0d", X"7d", X"3c", X"74", X"99", 
    X"5d", X"b4", X"18", X"05", X"75", X"99", X"63", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"7e", 
    X"3c", X"74", X"99", X"5e", X"b4", X"18", X"0d", X"7f", 
    X"3c", X"74", X"99", X"5f", X"b4", X"18", X"05", X"75", 
    X"99", X"64", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"74", X"99", X"54", X"3c", X"f5", X"e0", 
    X"b4", X"18", X"05", X"75", X"99", X"65", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"60", 
    X"99", X"53", X"60", X"3c", X"85", X"60", X"e0", X"b4", 
    X"18", X"11", X"75", X"f0", X"99", X"53", X"f0", X"3c", 
    X"85", X"f0", X"e0", X"b4", X"18", X"05", X"75", X"99", 
    X"66", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"60", X"3c", X"74", X"99", X"52", X"60", 
    X"e5", X"60", X"b4", X"18", X"05", X"75", X"99", X"67", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", X"99", 
    X"49", X"75", X"60", X"51", X"74", X"92", X"45", X"60", 
    X"b4", X"d3", X"29", X"78", X"60", X"76", X"51", X"74", 
    X"92", X"46", X"b4", X"d3", X"1f", X"79", X"31", X"77", 
    X"51", X"74", X"92", X"47", X"b4", X"d3", X"15", X"78", 
    X"51", X"74", X"92", X"48", X"b4", X"d3", X"0d", X"79", 
    X"51", X"74", X"92", X"49", X"b4", X"d3", X"05", X"75", 
    X"99", X"61", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"7a", X"51", X"74", X"92", X"4a", X"b4", 
    X"d3", X"0d", X"7b", X"51", X"74", X"92", X"4b", X"b4", 
    X"d3", X"05", X"75", X"99", X"62", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7c", X"51", X"74", 
    X"92", X"4c", X"b4", X"d3", X"0d", X"7d", X"51", X"74", 
    X"92", X"4d", X"b4", X"d3", X"05", X"75", X"99", X"63", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"7e", X"51", X"74", X"92", X"4e", X"b4", X"d3", X"0d", 
    X"7f", X"51", X"74", X"92", X"4f", X"b4", X"d3", X"05", 
    X"75", X"99", X"64", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"74", X"92", X"44", X"51", X"f5", 
    X"e0", X"b4", X"d3", X"05", X"75", X"99", X"65", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"60", X"92", X"43", X"60", X"51", X"85", X"60", X"e0", 
    X"b4", X"d3", X"11", X"75", X"f0", X"92", X"43", X"f0", 
    X"51", X"85", X"f0", X"e0", X"b4", X"d3", X"05", X"75", 
    X"99", X"66", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"60", X"51", X"74", X"92", X"42", 
    X"60", X"e5", X"60", X"b4", X"d3", X"05", X"75", X"99", 
    X"67", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", 
    X"99", X"4a", X"75", X"60", X"51", X"74", X"33", X"65", 
    X"60", X"b4", X"62", X"29", X"78", X"60", X"76", X"51", 
    X"74", X"33", X"66", X"b4", X"62", X"1f", X"79", X"31", 
    X"77", X"51", X"74", X"33", X"67", X"b4", X"62", X"15", 
    X"78", X"51", X"74", X"33", X"68", X"b4", X"62", X"0d", 
    X"79", X"51", X"74", X"33", X"69", X"b4", X"62", X"05", 
    X"75", X"99", X"61", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"7a", X"51", X"74", X"33", X"6a", 
    X"b4", X"62", X"0d", X"7b", X"51", X"74", X"33", X"6b", 
    X"b4", X"62", X"05", X"75", X"99", X"62", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7c", X"51", 
    X"74", X"33", X"6c", X"b4", X"62", X"0d", X"7d", X"51", 
    X"74", X"33", X"6d", X"b4", X"62", X"05", X"75", X"99", 
    X"63", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"7e", X"51", X"74", X"33", X"6e", X"b4", X"62", 
    X"0d", X"7f", X"51", X"74", X"33", X"6f", X"b4", X"62", 
    X"05", X"75", X"99", X"64", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"74", X"33", X"64", X"51", 
    X"f5", X"e0", X"b4", X"62", X"05", X"75", X"99", X"65", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"75", X"60", X"33", X"63", X"60", X"51", X"85", X"60", 
    X"e0", X"b4", X"62", X"11", X"75", X"f0", X"33", X"63", 
    X"f0", X"51", X"85", X"f0", X"e0", X"b4", X"62", X"05", 
    X"75", X"99", X"66", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"75", X"60", X"51", X"74", X"33", 
    X"62", X"60", X"e5", X"60", X"b4", X"62", X"05", X"75", 
    X"99", X"67", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"99", X"0d", X"75", X"99", X"0a", 
    X"75", X"99", X"4b", X"75", X"60", X"03", X"74", X"04", 
    X"14", X"60", X"19", X"d5", X"60", X"fa", X"b4", X"01", 
    X"13", X"75", X"f0", X"03", X"74", X"04", X"14", X"60", 
    X"0b", X"d5", X"f0", X"fa", X"b4", X"01", X"05", X"75", 
    X"99", X"61", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"78", X"03", X"74", X"04", X"14", X"60", 
    X"5e", X"d8", X"fb", X"b4", X"01", X"59", X"79", X"03", 
    X"74", X"04", X"14", X"60", X"52", X"d9", X"fb", X"b4", 
    X"01", X"4d", X"7a", X"03", X"74", X"04", X"14", X"60", 
    X"46", X"da", X"fb", X"b4", X"01", X"41", X"7b", X"03", 
    X"74", X"04", X"14", X"60", X"3a", X"db", X"fb", X"b4", 
    X"01", X"35", X"7c", X"03", X"74", X"04", X"14", X"60", 
    X"2e", X"dc", X"fb", X"b4", X"01", X"29", X"7d", X"03", 
    X"74", X"04", X"14", X"60", X"22", X"dd", X"fb", X"b4", 
    X"01", X"1d", X"7e", X"03", X"74", X"04", X"14", X"60", 
    X"16", X"de", X"fb", X"b4", X"01", X"11", X"7f", X"03", 
    X"74", X"04", X"14", X"60", X"0a", X"df", X"fb", X"b4", 
    X"01", X"05", X"75", X"99", X"62", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", X"0d", 
    X"75", X"99", X"0a", X"75", X"99", X"4c", X"75", X"99", 
    X"30", X"75", X"60", X"51", X"74", X"33", X"c3", X"25", 
    X"60", X"85", X"d0", X"70", X"b4", X"84", X"6b", X"e5", 
    X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", X"70", 
    X"61", X"78", X"60", X"76", X"51", X"74", X"33", X"c3", 
    X"26", X"85", X"d0", X"70", X"b4", X"84", X"53", X"e5", 
    X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", X"70", 
    X"49", X"79", X"31", X"77", X"51", X"74", X"33", X"c3", 
    X"27", X"85", X"d0", X"70", X"b4", X"84", X"3b", X"e5", 
    X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", X"70", 
    X"31", X"78", X"51", X"74", X"33", X"c3", X"28", X"85", 
    X"d0", X"70", X"b4", X"84", X"25", X"e5", X"70", X"54", 
    X"c4", X"64", X"04", X"54", X"fe", X"70", X"1b", X"79", 
    X"51", X"74", X"33", X"c3", X"29", X"85", X"d0", X"70", 
    X"b4", X"84", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"04", X"54", X"fe", X"70", X"05", X"75", X"99", X"61", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"7a", X"51", X"74", X"33", X"c3", X"2a", X"85", X"d0", 
    X"70", X"b4", X"84", X"25", X"e5", X"70", X"54", X"c4", 
    X"64", X"04", X"54", X"fe", X"70", X"1b", X"7b", X"51", 
    X"74", X"33", X"c3", X"2b", X"85", X"d0", X"70", X"b4", 
    X"84", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"04", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"62", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"7c", 
    X"51", X"74", X"33", X"c3", X"2c", X"85", X"d0", X"70", 
    X"b4", X"84", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"04", X"54", X"fe", X"70", X"1b", X"7d", X"51", X"74", 
    X"33", X"c3", X"2d", X"85", X"d0", X"70", X"b4", X"84", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"04", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"63", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7e", X"51", 
    X"74", X"33", X"c3", X"2e", X"85", X"d0", X"70", X"b4", 
    X"84", X"25", X"e5", X"70", X"54", X"c4", X"64", X"04", 
    X"54", X"fe", X"70", X"1b", X"7f", X"51", X"74", X"33", 
    X"c3", X"2f", X"85", X"d0", X"70", X"b4", X"84", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"64", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"74", X"33", X"c3", 
    X"24", X"51", X"85", X"d0", X"70", X"f5", X"e0", X"b4", 
    X"84", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"04", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"65", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"99", X"31", X"75", X"60", X"81", X"74", X"93", X"c3", 
    X"25", X"60", X"85", X"d0", X"70", X"b4", X"14", X"6b", 
    X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", X"fe", 
    X"70", X"61", X"78", X"60", X"76", X"81", X"74", X"93", 
    X"c3", X"26", X"85", X"d0", X"70", X"b4", X"14", X"53", 
    X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", X"fe", 
    X"70", X"49", X"79", X"31", X"77", X"81", X"74", X"93", 
    X"c3", X"27", X"85", X"d0", X"70", X"b4", X"14", X"3b", 
    X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", X"fe", 
    X"70", X"31", X"78", X"81", X"74", X"93", X"c3", X"28", 
    X"85", X"d0", X"70", X"b4", X"14", X"25", X"e5", X"70", 
    X"54", X"c4", X"64", X"84", X"54", X"fe", X"70", X"1b", 
    X"79", X"81", X"74", X"93", X"c3", X"29", X"85", X"d0", 
    X"70", X"b4", X"14", X"0f", X"e5", X"70", X"54", X"c4", 
    X"64", X"84", X"54", X"fe", X"70", X"05", X"75", X"99", 
    X"61", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"7a", X"81", X"74", X"93", X"c3", X"2a", X"85", 
    X"d0", X"70", X"b4", X"14", X"25", X"e5", X"70", X"54", 
    X"c4", X"64", X"84", X"54", X"fe", X"70", X"1b", X"7b", 
    X"81", X"74", X"93", X"c3", X"2b", X"85", X"d0", X"70", 
    X"b4", X"14", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"84", X"54", X"fe", X"70", X"05", X"75", X"99", X"62", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"7c", X"81", X"74", X"93", X"c3", X"2c", X"85", X"d0", 
    X"70", X"b4", X"14", X"25", X"e5", X"70", X"54", X"c4", 
    X"64", X"84", X"54", X"fe", X"70", X"1b", X"7d", X"81", 
    X"74", X"93", X"c3", X"2d", X"85", X"d0", X"70", X"b4", 
    X"14", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"84", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"63", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"7e", 
    X"81", X"74", X"93", X"c3", X"2e", X"85", X"d0", X"70", 
    X"b4", X"14", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"84", X"54", X"fe", X"70", X"1b", X"7f", X"81", X"74", 
    X"93", X"c3", X"2f", X"85", X"d0", X"70", X"b4", X"14", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"64", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"74", X"93", 
    X"c3", X"24", X"81", X"85", X"d0", X"70", X"f5", X"e0", 
    X"b4", X"14", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"84", X"54", X"fe", X"70", X"05", X"75", X"99", X"65", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"75", X"99", X"32", X"75", X"60", X"88", X"74", X"98", 
    X"c3", X"25", X"60", X"85", X"d0", X"70", X"b4", X"20", 
    X"6b", X"e5", X"70", X"54", X"c4", X"64", X"c4", X"54", 
    X"fe", X"70", X"61", X"78", X"60", X"76", X"88", X"74", 
    X"98", X"c3", X"26", X"85", X"d0", X"70", X"b4", X"20", 
    X"53", X"e5", X"70", X"54", X"c4", X"64", X"c4", X"54", 
    X"fe", X"70", X"49", X"79", X"31", X"77", X"88", X"74", 
    X"98", X"c3", X"27", X"85", X"d0", X"70", X"b4", X"20", 
    X"3b", X"e5", X"70", X"54", X"c4", X"64", X"c4", X"54", 
    X"fe", X"70", X"31", X"78", X"88", X"74", X"98", X"c3", 
    X"28", X"85", X"d0", X"70", X"b4", X"20", X"25", X"e5", 
    X"70", X"54", X"c4", X"64", X"c4", X"54", X"fe", X"70", 
    X"1b", X"79", X"88", X"74", X"98", X"c3", X"29", X"85", 
    X"d0", X"70", X"b4", X"20", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"c4", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"61", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"7a", X"88", X"74", X"98", X"c3", X"2a", 
    X"85", X"d0", X"70", X"b4", X"20", X"25", X"e5", X"70", 
    X"54", X"c4", X"64", X"c4", X"54", X"fe", X"70", X"1b", 
    X"7b", X"88", X"74", X"98", X"c3", X"2b", X"85", X"d0", 
    X"70", X"b4", X"20", X"0f", X"e5", X"70", X"54", X"c4", 
    X"64", X"c4", X"54", X"fe", X"70", X"05", X"75", X"99", 
    X"62", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"7c", X"88", X"74", X"98", X"c3", X"2c", X"85", 
    X"d0", X"70", X"b4", X"20", X"25", X"e5", X"70", X"54", 
    X"c4", X"64", X"c4", X"54", X"fe", X"70", X"1b", X"7d", 
    X"88", X"74", X"98", X"c3", X"2d", X"85", X"d0", X"70", 
    X"b4", X"20", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"c4", X"54", X"fe", X"70", X"05", X"75", X"99", X"63", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"7e", X"88", X"74", X"98", X"c3", X"2e", X"85", X"d0", 
    X"70", X"b4", X"20", X"25", X"e5", X"70", X"54", X"c4", 
    X"64", X"c4", X"54", X"fe", X"70", X"1b", X"7f", X"88", 
    X"74", X"98", X"c3", X"2f", X"85", X"d0", X"70", X"b4", 
    X"20", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c4", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"64", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"74", 
    X"98", X"c3", X"24", X"88", X"85", X"d0", X"70", X"f5", 
    X"e0", X"b4", X"20", X"0f", X"e5", X"70", X"54", X"c4", 
    X"64", X"c4", X"54", X"fe", X"70", X"05", X"75", X"99", 
    X"65", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"75", X"99", X"33", X"75", X"60", X"43", X"74", 
    X"fb", X"c3", X"25", X"60", X"85", X"d0", X"70", X"b4", 
    X"3e", X"6b", X"e5", X"70", X"54", X"c4", X"64", X"80", 
    X"54", X"fe", X"70", X"61", X"78", X"60", X"76", X"43", 
    X"74", X"fb", X"c3", X"26", X"85", X"d0", X"70", X"b4", 
    X"3e", X"53", X"e5", X"70", X"54", X"c4", X"64", X"80", 
    X"54", X"fe", X"70", X"49", X"79", X"31", X"77", X"43", 
    X"74", X"fb", X"c3", X"27", X"85", X"d0", X"70", X"b4", 
    X"3e", X"3b", X"e5", X"70", X"54", X"c4", X"64", X"80", 
    X"54", X"fe", X"70", X"31", X"78", X"43", X"74", X"fb", 
    X"c3", X"28", X"85", X"d0", X"70", X"b4", X"3e", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"80", X"54", X"fe", 
    X"70", X"1b", X"79", X"43", X"74", X"fb", X"c3", X"29", 
    X"85", X"d0", X"70", X"b4", X"3e", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"80", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"61", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"7a", X"43", X"74", X"fb", X"c3", 
    X"2a", X"85", X"d0", X"70", X"b4", X"3e", X"25", X"e5", 
    X"70", X"54", X"c4", X"64", X"80", X"54", X"fe", X"70", 
    X"1b", X"7b", X"43", X"74", X"fb", X"c3", X"2b", X"85", 
    X"d0", X"70", X"b4", X"3e", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"80", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"62", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"7c", X"43", X"74", X"fb", X"c3", X"2c", 
    X"85", X"d0", X"70", X"b4", X"3e", X"25", X"e5", X"70", 
    X"54", X"c4", X"64", X"80", X"54", X"fe", X"70", X"1b", 
    X"7d", X"43", X"74", X"fb", X"c3", X"2d", X"85", X"d0", 
    X"70", X"b4", X"3e", X"0f", X"e5", X"70", X"54", X"c4", 
    X"64", X"80", X"54", X"fe", X"70", X"05", X"75", X"99", 
    X"63", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"7e", X"43", X"74", X"fb", X"c3", X"2e", X"85", 
    X"d0", X"70", X"b4", X"3e", X"25", X"e5", X"70", X"54", 
    X"c4", X"64", X"80", X"54", X"fe", X"70", X"1b", X"7f", 
    X"43", X"74", X"fb", X"c3", X"2f", X"85", X"d0", X"70", 
    X"b4", X"3e", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"80", X"54", X"fe", X"70", X"05", X"75", X"99", X"64", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"74", X"fb", X"c3", X"24", X"43", X"85", X"d0", X"70", 
    X"f5", X"e0", X"b4", X"3e", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"80", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"65", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"99", X"0d", X"75", X"99", X"0a", 
    X"75", X"99", X"4d", X"75", X"99", X"30", X"75", X"60", 
    X"51", X"74", X"33", X"c3", X"35", X"60", X"85", X"d0", 
    X"70", X"b4", X"84", X"6b", X"e5", X"70", X"54", X"c4", 
    X"64", X"04", X"54", X"fe", X"70", X"61", X"78", X"60", 
    X"76", X"51", X"74", X"33", X"c3", X"36", X"85", X"d0", 
    X"70", X"b4", X"84", X"53", X"e5", X"70", X"54", X"c4", 
    X"64", X"04", X"54", X"fe", X"70", X"49", X"79", X"31", 
    X"77", X"51", X"74", X"33", X"c3", X"37", X"85", X"d0", 
    X"70", X"b4", X"84", X"3b", X"e5", X"70", X"54", X"c4", 
    X"64", X"04", X"54", X"fe", X"70", X"31", X"78", X"51", 
    X"74", X"33", X"c3", X"38", X"85", X"d0", X"70", X"b4", 
    X"84", X"25", X"e5", X"70", X"54", X"c4", X"64", X"04", 
    X"54", X"fe", X"70", X"1b", X"79", X"51", X"74", X"33", 
    X"c3", X"39", X"85", X"d0", X"70", X"b4", X"84", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"61", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7a", X"51", X"74", 
    X"33", X"c3", X"3a", X"85", X"d0", X"70", X"b4", X"84", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"04", X"54", 
    X"fe", X"70", X"1b", X"7b", X"51", X"74", X"33", X"c3", 
    X"3b", X"85", X"d0", X"70", X"b4", X"84", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"62", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7c", X"51", X"74", X"33", 
    X"c3", X"3c", X"85", X"d0", X"70", X"b4", X"84", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", 
    X"70", X"1b", X"7d", X"51", X"74", X"33", X"c3", X"3d", 
    X"85", X"d0", X"70", X"b4", X"84", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"04", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"63", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"7e", X"51", X"74", X"33", X"c3", 
    X"3e", X"85", X"d0", X"70", X"b4", X"84", X"25", X"e5", 
    X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", X"70", 
    X"1b", X"7f", X"51", X"74", X"33", X"c3", X"3f", X"85", 
    X"d0", X"70", X"b4", X"84", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"04", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"64", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"74", X"33", X"c3", X"34", X"51", X"85", 
    X"d0", X"70", X"f5", X"e0", X"b4", X"84", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"04", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"65", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"99", X"31", X"75", 
    X"60", X"81", X"74", X"93", X"c3", X"35", X"60", X"85", 
    X"d0", X"70", X"b4", X"14", X"6b", X"e5", X"70", X"54", 
    X"c4", X"64", X"84", X"54", X"fe", X"70", X"61", X"78", 
    X"60", X"76", X"81", X"74", X"93", X"c3", X"36", X"85", 
    X"d0", X"70", X"b4", X"14", X"53", X"e5", X"70", X"54", 
    X"c4", X"64", X"84", X"54", X"fe", X"70", X"49", X"79", 
    X"31", X"77", X"81", X"74", X"93", X"c3", X"37", X"85", 
    X"d0", X"70", X"b4", X"14", X"3b", X"e5", X"70", X"54", 
    X"c4", X"64", X"84", X"54", X"fe", X"70", X"31", X"78", 
    X"81", X"74", X"93", X"c3", X"38", X"85", X"d0", X"70", 
    X"b4", X"14", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"84", X"54", X"fe", X"70", X"1b", X"79", X"81", X"74", 
    X"93", X"c3", X"39", X"85", X"d0", X"70", X"b4", X"14", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"61", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7a", X"81", 
    X"74", X"93", X"c3", X"3a", X"85", X"d0", X"70", X"b4", 
    X"14", X"25", X"e5", X"70", X"54", X"c4", X"64", X"84", 
    X"54", X"fe", X"70", X"1b", X"7b", X"81", X"74", X"93", 
    X"c3", X"3b", X"85", X"d0", X"70", X"b4", X"14", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"62", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7c", X"81", X"74", 
    X"93", X"c3", X"3c", X"85", X"d0", X"70", X"b4", X"14", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", 
    X"fe", X"70", X"1b", X"7d", X"81", X"74", X"93", X"c3", 
    X"3d", X"85", X"d0", X"70", X"b4", X"14", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"84", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"63", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7e", X"81", X"74", X"93", 
    X"c3", X"3e", X"85", X"d0", X"70", X"b4", X"14", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", X"fe", 
    X"70", X"1b", X"7f", X"81", X"74", X"93", X"c3", X"3f", 
    X"85", X"d0", X"70", X"b4", X"14", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"84", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"64", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"74", X"93", X"c3", X"34", X"81", 
    X"85", X"d0", X"70", X"f5", X"e0", X"b4", X"14", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"84", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"65", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", X"32", 
    X"75", X"60", X"88", X"74", X"98", X"c3", X"35", X"60", 
    X"85", X"d0", X"70", X"b4", X"20", X"6b", X"e5", X"70", 
    X"54", X"c4", X"64", X"c4", X"54", X"fe", X"70", X"61", 
    X"78", X"60", X"76", X"88", X"74", X"98", X"c3", X"36", 
    X"85", X"d0", X"70", X"b4", X"20", X"53", X"e5", X"70", 
    X"54", X"c4", X"64", X"c4", X"54", X"fe", X"70", X"49", 
    X"79", X"31", X"77", X"88", X"74", X"98", X"c3", X"37", 
    X"85", X"d0", X"70", X"b4", X"20", X"3b", X"e5", X"70", 
    X"54", X"c4", X"64", X"c4", X"54", X"fe", X"70", X"31", 
    X"78", X"88", X"74", X"98", X"c3", X"38", X"85", X"d0", 
    X"70", X"b4", X"20", X"25", X"e5", X"70", X"54", X"c4", 
    X"64", X"c4", X"54", X"fe", X"70", X"1b", X"79", X"88", 
    X"74", X"98", X"c3", X"39", X"85", X"d0", X"70", X"b4", 
    X"20", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c4", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"61", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"7a", 
    X"88", X"74", X"98", X"c3", X"3a", X"85", X"d0", X"70", 
    X"b4", X"20", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"c4", X"54", X"fe", X"70", X"1b", X"7b", X"88", X"74", 
    X"98", X"c3", X"3b", X"85", X"d0", X"70", X"b4", X"20", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c4", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"62", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7c", X"88", 
    X"74", X"98", X"c3", X"3c", X"85", X"d0", X"70", X"b4", 
    X"20", X"25", X"e5", X"70", X"54", X"c4", X"64", X"c4", 
    X"54", X"fe", X"70", X"1b", X"7d", X"88", X"74", X"98", 
    X"c3", X"3d", X"85", X"d0", X"70", X"b4", X"20", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"c4", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"63", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7e", X"88", X"74", 
    X"98", X"c3", X"3e", X"85", X"d0", X"70", X"b4", X"20", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"c4", X"54", 
    X"fe", X"70", X"1b", X"7f", X"88", X"74", X"98", X"c3", 
    X"3f", X"85", X"d0", X"70", X"b4", X"20", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"c4", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"64", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"74", X"98", X"c3", X"34", 
    X"88", X"85", X"d0", X"70", X"f5", X"e0", X"b4", X"20", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c4", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"65", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", 
    X"33", X"75", X"60", X"88", X"74", X"98", X"d3", X"35", 
    X"60", X"85", X"d0", X"70", X"b4", X"21", X"6b", X"e5", 
    X"70", X"54", X"c4", X"64", X"c5", X"54", X"fe", X"70", 
    X"61", X"78", X"60", X"76", X"88", X"74", X"98", X"d3", 
    X"36", X"85", X"d0", X"70", X"b4", X"21", X"53", X"e5", 
    X"70", X"54", X"c4", X"64", X"c5", X"54", X"fe", X"70", 
    X"49", X"79", X"31", X"77", X"88", X"74", X"98", X"d3", 
    X"37", X"85", X"d0", X"70", X"b4", X"21", X"3b", X"e5", 
    X"70", X"54", X"c4", X"64", X"c5", X"54", X"fe", X"70", 
    X"31", X"78", X"88", X"74", X"98", X"d3", X"38", X"85", 
    X"d0", X"70", X"b4", X"21", X"25", X"e5", X"70", X"54", 
    X"c4", X"64", X"c5", X"54", X"fe", X"70", X"1b", X"79", 
    X"88", X"74", X"98", X"d3", X"39", X"85", X"d0", X"70", 
    X"b4", X"21", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"c5", X"54", X"fe", X"70", X"05", X"75", X"99", X"61", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"7a", X"88", X"74", X"98", X"d3", X"3a", X"85", X"d0", 
    X"70", X"b4", X"21", X"25", X"e5", X"70", X"54", X"c4", 
    X"64", X"c5", X"54", X"fe", X"70", X"1b", X"7b", X"88", 
    X"74", X"98", X"d3", X"3b", X"85", X"d0", X"70", X"b4", 
    X"21", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c5", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"62", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"7c", 
    X"88", X"74", X"98", X"d3", X"3c", X"85", X"d0", X"70", 
    X"b4", X"21", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"c5", X"54", X"fe", X"70", X"1b", X"7d", X"88", X"74", 
    X"98", X"d3", X"3d", X"85", X"d0", X"70", X"b4", X"21", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c5", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"63", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7e", X"88", 
    X"74", X"98", X"d3", X"3e", X"85", X"d0", X"70", X"b4", 
    X"21", X"25", X"e5", X"70", X"54", X"c4", X"64", X"c5", 
    X"54", X"fe", X"70", X"1b", X"7f", X"88", X"74", X"98", 
    X"d3", X"3f", X"85", X"d0", X"70", X"b4", X"21", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"c5", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"64", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"74", X"98", X"d3", 
    X"34", X"88", X"85", X"d0", X"70", X"f5", X"e0", X"b4", 
    X"21", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c5", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"65", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"99", X"34", X"75", X"60", X"43", X"74", X"fb", X"d3", 
    X"35", X"60", X"85", X"d0", X"70", X"b4", X"3f", X"6b", 
    X"e5", X"70", X"54", X"c4", X"64", X"81", X"54", X"fe", 
    X"70", X"61", X"78", X"60", X"76", X"43", X"74", X"fb", 
    X"d3", X"36", X"85", X"d0", X"70", X"b4", X"3f", X"53", 
    X"e5", X"70", X"54", X"c4", X"64", X"81", X"54", X"fe", 
    X"70", X"49", X"79", X"31", X"77", X"43", X"74", X"fb", 
    X"d3", X"37", X"85", X"d0", X"70", X"b4", X"3f", X"3b", 
    X"e5", X"70", X"54", X"c4", X"64", X"81", X"54", X"fe", 
    X"70", X"31", X"78", X"43", X"74", X"fb", X"d3", X"38", 
    X"85", X"d0", X"70", X"b4", X"3f", X"25", X"e5", X"70", 
    X"54", X"c4", X"64", X"81", X"54", X"fe", X"70", X"1b", 
    X"79", X"43", X"74", X"fb", X"d3", X"39", X"85", X"d0", 
    X"70", X"b4", X"3f", X"0f", X"e5", X"70", X"54", X"c4", 
    X"64", X"81", X"54", X"fe", X"70", X"05", X"75", X"99", 
    X"61", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"7a", X"43", X"74", X"fb", X"d3", X"3a", X"85", 
    X"d0", X"70", X"b4", X"3f", X"25", X"e5", X"70", X"54", 
    X"c4", X"64", X"81", X"54", X"fe", X"70", X"1b", X"7b", 
    X"43", X"74", X"fb", X"d3", X"3b", X"85", X"d0", X"70", 
    X"b4", X"3f", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"81", X"54", X"fe", X"70", X"05", X"75", X"99", X"62", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"7c", X"43", X"74", X"fb", X"d3", X"3c", X"85", X"d0", 
    X"70", X"b4", X"3f", X"25", X"e5", X"70", X"54", X"c4", 
    X"64", X"81", X"54", X"fe", X"70", X"1b", X"7d", X"43", 
    X"74", X"fb", X"d3", X"3d", X"85", X"d0", X"70", X"b4", 
    X"3f", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"81", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"63", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"7e", 
    X"43", X"74", X"fb", X"d3", X"3e", X"85", X"d0", X"70", 
    X"b4", X"3f", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"81", X"54", X"fe", X"70", X"1b", X"7f", X"43", X"74", 
    X"fb", X"d3", X"3f", X"85", X"d0", X"70", X"b4", X"3f", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"81", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"64", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"74", X"fb", 
    X"d3", X"34", X"43", X"85", X"d0", X"70", X"f5", X"e0", 
    X"b4", X"3f", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"81", X"54", X"fe", X"70", X"05", X"75", X"99", X"65", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", X"99", 
    X"4e", X"75", X"99", X"30", X"75", X"60", X"70", X"74", 
    X"73", X"c3", X"95", X"60", X"85", X"d0", X"70", X"b4", 
    X"03", X"6b", X"e5", X"70", X"54", X"c4", X"64", X"00", 
    X"54", X"fe", X"70", X"61", X"78", X"60", X"76", X"70", 
    X"74", X"73", X"c3", X"96", X"85", X"d0", X"70", X"b4", 
    X"03", X"53", X"e5", X"70", X"54", X"c4", X"64", X"00", 
    X"54", X"fe", X"70", X"49", X"79", X"31", X"77", X"70", 
    X"74", X"73", X"c3", X"97", X"85", X"d0", X"70", X"b4", 
    X"03", X"3b", X"e5", X"70", X"54", X"c4", X"64", X"00", 
    X"54", X"fe", X"70", X"31", X"78", X"70", X"74", X"73", 
    X"c3", X"98", X"85", X"d0", X"70", X"b4", X"03", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"00", X"54", X"fe", 
    X"70", X"1b", X"79", X"70", X"74", X"73", X"c3", X"99", 
    X"85", X"d0", X"70", X"b4", X"03", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"00", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"61", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"7a", X"70", X"74", X"73", X"c3", 
    X"9a", X"85", X"d0", X"70", X"b4", X"03", X"25", X"e5", 
    X"70", X"54", X"c4", X"64", X"00", X"54", X"fe", X"70", 
    X"1b", X"7b", X"70", X"74", X"73", X"c3", X"9b", X"85", 
    X"d0", X"70", X"b4", X"03", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"00", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"62", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"7c", X"70", X"74", X"73", X"c3", X"9c", 
    X"85", X"d0", X"70", X"b4", X"03", X"25", X"e5", X"70", 
    X"54", X"c4", X"64", X"00", X"54", X"fe", X"70", X"1b", 
    X"7d", X"70", X"74", X"73", X"c3", X"9d", X"85", X"d0", 
    X"70", X"b4", X"03", X"0f", X"e5", X"70", X"54", X"c4", 
    X"64", X"00", X"54", X"fe", X"70", X"05", X"75", X"99", 
    X"63", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"7e", X"70", X"74", X"73", X"c3", X"9e", X"85", 
    X"d0", X"70", X"b4", X"03", X"25", X"e5", X"70", X"54", 
    X"c4", X"64", X"00", X"54", X"fe", X"70", X"1b", X"7f", 
    X"70", X"74", X"73", X"c3", X"9f", X"85", X"d0", X"70", 
    X"b4", X"03", X"0f", X"e5", X"70", X"54", X"c4", X"64", 
    X"00", X"54", X"fe", X"70", X"05", X"75", X"99", X"64", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"74", X"73", X"c3", X"94", X"70", X"85", X"d0", X"70", 
    X"f5", X"e0", X"b4", X"03", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"00", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"65", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"99", X"31", X"75", X"60", X"70", 
    X"74", X"73", X"d3", X"95", X"60", X"85", X"d0", X"70", 
    X"b4", X"02", X"6b", X"e5", X"70", X"54", X"c4", X"64", 
    X"01", X"54", X"fe", X"70", X"61", X"78", X"60", X"76", 
    X"70", X"74", X"73", X"d3", X"96", X"85", X"d0", X"70", 
    X"b4", X"02", X"53", X"e5", X"70", X"54", X"c4", X"64", 
    X"01", X"54", X"fe", X"70", X"49", X"79", X"31", X"77", 
    X"70", X"74", X"73", X"d3", X"97", X"85", X"d0", X"70", 
    X"b4", X"02", X"3b", X"e5", X"70", X"54", X"c4", X"64", 
    X"01", X"54", X"fe", X"70", X"31", X"78", X"70", X"74", 
    X"73", X"d3", X"98", X"85", X"d0", X"70", X"b4", X"02", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"01", X"54", 
    X"fe", X"70", X"1b", X"79", X"70", X"74", X"73", X"d3", 
    X"99", X"85", X"d0", X"70", X"b4", X"02", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"01", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"61", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7a", X"70", X"74", X"73", 
    X"d3", X"9a", X"85", X"d0", X"70", X"b4", X"02", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"01", X"54", X"fe", 
    X"70", X"1b", X"7b", X"70", X"74", X"73", X"d3", X"9b", 
    X"85", X"d0", X"70", X"b4", X"02", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"01", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"62", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"7c", X"70", X"74", X"73", X"d3", 
    X"9c", X"85", X"d0", X"70", X"b4", X"02", X"25", X"e5", 
    X"70", X"54", X"c4", X"64", X"01", X"54", X"fe", X"70", 
    X"1b", X"7d", X"70", X"74", X"73", X"d3", X"9d", X"85", 
    X"d0", X"70", X"b4", X"02", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"01", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"63", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"7e", X"70", X"74", X"73", X"d3", X"9e", 
    X"85", X"d0", X"70", X"b4", X"02", X"25", X"e5", X"70", 
    X"54", X"c4", X"64", X"01", X"54", X"fe", X"70", X"1b", 
    X"7f", X"70", X"74", X"73", X"d3", X"9f", X"85", X"d0", 
    X"70", X"b4", X"02", X"0f", X"e5", X"70", X"54", X"c4", 
    X"64", X"01", X"54", X"fe", X"70", X"05", X"75", X"99", 
    X"64", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"74", X"73", X"d3", X"94", X"70", X"85", X"d0", 
    X"70", X"f5", X"e0", X"b4", X"02", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"01", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"65", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"75", X"99", X"32", X"75", X"60", 
    X"c3", X"74", X"c5", X"c3", X"95", X"60", X"85", X"d0", 
    X"70", X"b4", X"02", X"6b", X"e5", X"70", X"54", X"c4", 
    X"64", X"00", X"54", X"fe", X"70", X"61", X"78", X"60", 
    X"76", X"c3", X"74", X"c5", X"c3", X"96", X"85", X"d0", 
    X"70", X"b4", X"02", X"53", X"e5", X"70", X"54", X"c4", 
    X"64", X"00", X"54", X"fe", X"70", X"49", X"79", X"31", 
    X"77", X"c3", X"74", X"c5", X"c3", X"97", X"85", X"d0", 
    X"70", X"b4", X"02", X"3b", X"e5", X"70", X"54", X"c4", 
    X"64", X"00", X"54", X"fe", X"70", X"31", X"78", X"c3", 
    X"74", X"c5", X"c3", X"98", X"85", X"d0", X"70", X"b4", 
    X"02", X"25", X"e5", X"70", X"54", X"c4", X"64", X"00", 
    X"54", X"fe", X"70", X"1b", X"79", X"c3", X"74", X"c5", 
    X"c3", X"99", X"85", X"d0", X"70", X"b4", X"02", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"00", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"61", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7a", X"c3", X"74", 
    X"c5", X"c3", X"9a", X"85", X"d0", X"70", X"b4", X"02", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"00", X"54", 
    X"fe", X"70", X"1b", X"7b", X"c3", X"74", X"c5", X"c3", 
    X"9b", X"85", X"d0", X"70", X"b4", X"02", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"00", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"62", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7c", X"c3", X"74", X"c5", 
    X"c3", X"9c", X"85", X"d0", X"70", X"b4", X"02", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"00", X"54", X"fe", 
    X"70", X"1b", X"7d", X"c3", X"74", X"c5", X"c3", X"9d", 
    X"85", X"d0", X"70", X"b4", X"02", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"00", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"63", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"7e", X"c3", X"74", X"c5", X"c3", 
    X"9e", X"85", X"d0", X"70", X"b4", X"02", X"25", X"e5", 
    X"70", X"54", X"c4", X"64", X"00", X"54", X"fe", X"70", 
    X"1b", X"7f", X"c3", X"74", X"c5", X"c3", X"9f", X"85", 
    X"d0", X"70", X"b4", X"02", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"00", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"64", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"74", X"c5", X"c3", X"94", X"c3", X"85", 
    X"d0", X"70", X"f5", X"e0", X"b4", X"02", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"00", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"65", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"99", X"33", X"75", 
    X"60", X"c3", X"74", X"c5", X"d3", X"95", X"60", X"85", 
    X"d0", X"70", X"b4", X"01", X"6b", X"e5", X"70", X"54", 
    X"c4", X"64", X"01", X"54", X"fe", X"70", X"61", X"78", 
    X"60", X"76", X"c3", X"74", X"c5", X"d3", X"96", X"85", 
    X"d0", X"70", X"b4", X"01", X"53", X"e5", X"70", X"54", 
    X"c4", X"64", X"01", X"54", X"fe", X"70", X"49", X"79", 
    X"31", X"77", X"c3", X"74", X"c5", X"d3", X"97", X"85", 
    X"d0", X"70", X"b4", X"01", X"3b", X"e5", X"70", X"54", 
    X"c4", X"64", X"01", X"54", X"fe", X"70", X"31", X"78", 
    X"c3", X"74", X"c5", X"d3", X"98", X"85", X"d0", X"70", 
    X"b4", X"01", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"01", X"54", X"fe", X"70", X"1b", X"79", X"c3", X"74", 
    X"c5", X"d3", X"99", X"85", X"d0", X"70", X"b4", X"01", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"01", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"61", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7a", X"c3", 
    X"74", X"c5", X"d3", X"9a", X"85", X"d0", X"70", X"b4", 
    X"01", X"25", X"e5", X"70", X"54", X"c4", X"64", X"01", 
    X"54", X"fe", X"70", X"1b", X"7b", X"c3", X"74", X"c5", 
    X"d3", X"9b", X"85", X"d0", X"70", X"b4", X"01", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"01", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"62", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7c", X"c3", X"74", 
    X"c5", X"d3", X"9c", X"85", X"d0", X"70", X"b4", X"01", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"01", X"54", 
    X"fe", X"70", X"1b", X"7d", X"c3", X"74", X"c5", X"d3", 
    X"9d", X"85", X"d0", X"70", X"b4", X"01", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"01", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"63", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7e", X"c3", X"74", X"c5", 
    X"d3", X"9e", X"85", X"d0", X"70", X"b4", X"01", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"01", X"54", X"fe", 
    X"70", X"1b", X"7f", X"c3", X"74", X"c5", X"d3", X"9f", 
    X"85", X"d0", X"70", X"b4", X"01", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"01", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"64", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"74", X"c5", X"d3", X"94", X"c3", 
    X"85", X"d0", X"70", X"f5", X"e0", X"b4", X"01", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"01", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"65", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", X"34", 
    X"75", X"60", X"01", X"74", X"00", X"c3", X"95", X"60", 
    X"85", X"d0", X"70", X"b4", X"ff", X"6b", X"e5", X"70", 
    X"54", X"c4", X"64", X"c0", X"54", X"fe", X"70", X"61", 
    X"78", X"60", X"76", X"01", X"74", X"00", X"c3", X"96", 
    X"85", X"d0", X"70", X"b4", X"ff", X"53", X"e5", X"70", 
    X"54", X"c4", X"64", X"c0", X"54", X"fe", X"70", X"49", 
    X"79", X"31", X"77", X"01", X"74", X"00", X"c3", X"97", 
    X"85", X"d0", X"70", X"b4", X"ff", X"3b", X"e5", X"70", 
    X"54", X"c4", X"64", X"c0", X"54", X"fe", X"70", X"31", 
    X"78", X"01", X"74", X"00", X"c3", X"98", X"85", X"d0", 
    X"70", X"b4", X"ff", X"25", X"e5", X"70", X"54", X"c4", 
    X"64", X"c0", X"54", X"fe", X"70", X"1b", X"79", X"01", 
    X"74", X"00", X"c3", X"99", X"85", X"d0", X"70", X"b4", 
    X"ff", X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c0", 
    X"54", X"fe", X"70", X"05", X"75", X"99", X"61", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"7a", 
    X"01", X"74", X"00", X"c3", X"9a", X"85", X"d0", X"70", 
    X"b4", X"ff", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"c0", X"54", X"fe", X"70", X"1b", X"7b", X"01", X"74", 
    X"00", X"c3", X"9b", X"85", X"d0", X"70", X"b4", X"ff", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"c0", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"62", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7c", X"01", 
    X"74", X"00", X"c3", X"9c", X"85", X"d0", X"70", X"b4", 
    X"ff", X"25", X"e5", X"70", X"54", X"c4", X"64", X"c0", 
    X"54", X"fe", X"70", X"1b", X"7d", X"01", X"74", X"00", 
    X"c3", X"9d", X"85", X"d0", X"70", X"b4", X"ff", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"c0", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"63", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7e", X"01", X"74", 
    X"00", X"c3", X"9e", X"85", X"d0", X"70", X"b4", X"ff", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"c0", X"54", 
    X"fe", X"70", X"1b", X"7f", X"01", X"74", X"00", X"c3", 
    X"9f", X"85", X"d0", X"70", X"b4", X"ff", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"c0", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"64", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"99", X"35", X"75", 
    X"60", X"10", X"74", X"0a", X"c3", X"95", X"60", X"85", 
    X"d0", X"70", X"b4", X"fa", X"6b", X"e5", X"70", X"54", 
    X"c4", X"64", X"80", X"54", X"fe", X"70", X"61", X"78", 
    X"60", X"76", X"10", X"74", X"0a", X"c3", X"96", X"85", 
    X"d0", X"70", X"b4", X"fa", X"53", X"e5", X"70", X"54", 
    X"c4", X"64", X"80", X"54", X"fe", X"70", X"49", X"79", 
    X"31", X"77", X"10", X"74", X"0a", X"c3", X"97", X"85", 
    X"d0", X"70", X"b4", X"fa", X"3b", X"e5", X"70", X"54", 
    X"c4", X"64", X"80", X"54", X"fe", X"70", X"31", X"78", 
    X"10", X"74", X"0a", X"c3", X"98", X"85", X"d0", X"70", 
    X"b4", X"fa", X"25", X"e5", X"70", X"54", X"c4", X"64", 
    X"80", X"54", X"fe", X"70", X"1b", X"79", X"10", X"74", 
    X"0a", X"c3", X"99", X"85", X"d0", X"70", X"b4", X"fa", 
    X"0f", X"e5", X"70", X"54", X"c4", X"64", X"80", X"54", 
    X"fe", X"70", X"05", X"75", X"99", X"61", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"7a", X"10", 
    X"74", X"0a", X"c3", X"9a", X"85", X"d0", X"70", X"b4", 
    X"fa", X"25", X"e5", X"70", X"54", X"c4", X"64", X"80", 
    X"54", X"fe", X"70", X"1b", X"7b", X"10", X"74", X"0a", 
    X"c3", X"9b", X"85", X"d0", X"70", X"b4", X"fa", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"80", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"62", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7c", X"10", X"74", 
    X"0a", X"c3", X"9c", X"85", X"d0", X"70", X"b4", X"fa", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"80", X"54", 
    X"fe", X"70", X"1b", X"7d", X"10", X"74", X"0a", X"c3", 
    X"9d", X"85", X"d0", X"70", X"b4", X"fa", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"80", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"63", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7e", X"10", X"74", X"0a", 
    X"c3", X"9e", X"85", X"d0", X"70", X"b4", X"fa", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"80", X"54", X"fe", 
    X"70", X"1b", X"7f", X"10", X"74", X"0a", X"c3", X"9f", 
    X"85", X"d0", X"70", X"b4", X"fa", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"80", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"64", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"75", X"99", X"36", X"75", X"60", 
    X"10", X"74", X"0a", X"d3", X"95", X"60", X"85", X"d0", 
    X"70", X"b4", X"f9", X"6b", X"e5", X"70", X"54", X"c4", 
    X"64", X"81", X"54", X"fe", X"70", X"61", X"78", X"60", 
    X"76", X"10", X"74", X"0a", X"d3", X"96", X"85", X"d0", 
    X"70", X"b4", X"f9", X"53", X"e5", X"70", X"54", X"c4", 
    X"64", X"81", X"54", X"fe", X"70", X"49", X"79", X"31", 
    X"77", X"10", X"74", X"0a", X"d3", X"97", X"85", X"d0", 
    X"70", X"b4", X"f9", X"3b", X"e5", X"70", X"54", X"c4", 
    X"64", X"81", X"54", X"fe", X"70", X"31", X"78", X"10", 
    X"74", X"0a", X"d3", X"98", X"85", X"d0", X"70", X"b4", 
    X"f9", X"25", X"e5", X"70", X"54", X"c4", X"64", X"81", 
    X"54", X"fe", X"70", X"1b", X"79", X"10", X"74", X"0a", 
    X"d3", X"99", X"85", X"d0", X"70", X"b4", X"f9", X"0f", 
    X"e5", X"70", X"54", X"c4", X"64", X"81", X"54", X"fe", 
    X"70", X"05", X"75", X"99", X"61", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"7a", X"10", X"74", 
    X"0a", X"d3", X"9a", X"85", X"d0", X"70", X"b4", X"f9", 
    X"25", X"e5", X"70", X"54", X"c4", X"64", X"81", X"54", 
    X"fe", X"70", X"1b", X"7b", X"10", X"74", X"0a", X"d3", 
    X"9b", X"85", X"d0", X"70", X"b4", X"f9", X"0f", X"e5", 
    X"70", X"54", X"c4", X"64", X"81", X"54", X"fe", X"70", 
    X"05", X"75", X"99", X"62", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"7c", X"10", X"74", X"0a", 
    X"d3", X"9c", X"85", X"d0", X"70", X"b4", X"f9", X"25", 
    X"e5", X"70", X"54", X"c4", X"64", X"81", X"54", X"fe", 
    X"70", X"1b", X"7d", X"10", X"74", X"0a", X"d3", X"9d", 
    X"85", X"d0", X"70", X"b4", X"f9", X"0f", X"e5", X"70", 
    X"54", X"c4", X"64", X"81", X"54", X"fe", X"70", X"05", 
    X"75", X"99", X"63", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"7e", X"10", X"74", X"0a", X"d3", 
    X"9e", X"85", X"d0", X"70", X"b4", X"f9", X"25", X"e5", 
    X"70", X"54", X"c4", X"64", X"81", X"54", X"fe", X"70", 
    X"1b", X"7f", X"10", X"74", X"0a", X"d3", X"9f", X"85", 
    X"d0", X"70", X"b4", X"f9", X"0f", X"e5", X"70", X"54", 
    X"c4", X"64", X"81", X"54", X"fe", X"70", X"05", X"75", 
    X"99", X"64", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"99", X"0d", X"75", X"99", X"0a", 
    X"75", X"99", X"4f", X"75", X"81", X"9f", X"75", X"60", 
    X"12", X"78", X"a0", X"76", X"00", X"c0", X"60", X"e6", 
    X"b4", X"12", X"0a", X"e5", X"81", X"b4", X"a0", X"05", 
    X"75", X"99", X"61", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"75", X"61", X"00", X"e4", X"d0", 
    X"61", X"79", X"61", X"e7", X"b4", X"12", X"0a", X"e5", 
    X"81", X"b4", X"9f", X"05", X"75", X"99", X"62", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"81", X"9f", X"75", X"f0", X"42", X"78", X"a0", X"76", 
    X"00", X"c0", X"f0", X"e6", X"b4", X"42", X"0a", X"e5", 
    X"81", X"b4", X"a0", X"05", X"75", X"99", X"63", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"f0", X"00", X"e4", X"d0", X"f0", X"e5", X"f0", X"b4", 
    X"42", X"0a", X"e5", X"81", X"b4", X"9f", X"05", X"75", 
    X"99", X"64", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"75", X"99", X"0d", X"75", X"99", X"0a", 
    X"75", X"99", X"50", X"75", X"83", X"65", X"75", X"82", 
    X"43", X"90", X"01", X"23", X"e5", X"83", X"b4", X"01", 
    X"0a", X"e5", X"82", X"b4", X"23", X"05", X"75", X"99", 
    X"61", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"90", X"00", X"13", X"74", X"55", X"f0", X"a3", 
    X"f4", X"f0", X"90", X"00", X"13", X"e0", X"b4", X"55", 
    X"0a", X"a3", X"e0", X"b4", X"aa", X"05", X"75", X"99", 
    X"62", X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", 
    X"01", X"74", X"79", X"90", X"00", X"13", X"78", X"13", 
    X"79", X"14", X"f2", X"14", X"e0", X"b4", X"79", X"0d", 
    X"a3", X"74", X"97", X"f3", X"e0", X"b4", X"97", X"05", 
    X"75", X"99", X"63", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"74", X"79", X"90", X"00", X"13", 
    X"78", X"13", X"79", X"14", X"f0", X"14", X"e2", X"b4", 
    X"79", X"0e", X"74", X"97", X"a3", X"f0", X"14", X"e3", 
    X"b4", X"97", X"05", X"75", X"99", X"64", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", 
    X"0d", X"75", X"99", X"0a", X"75", X"99", X"51", X"74", 
    X"03", X"24", X"02", X"83", X"80", X"04", X"07", X"13", 
    X"19", X"21", X"b4", X"21", X"05", X"75", X"99", X"61", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"90", X"22", X"b6", X"74", X"00", X"93", X"b4", X"07", 
    X"17", X"74", X"01", X"93", X"b4", X"13", X"11", X"74", 
    X"02", X"93", X"b4", X"19", X"0b", X"74", X"03", X"93", 
    X"b4", X"21", X"05", X"75", X"99", X"62", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", 
    X"0d", X"75", X"99", X"0a", X"75", X"99", X"52", X"75", 
    X"81", X"4f", X"75", X"50", X"00", X"75", X"51", X"00", 
    X"75", X"52", X"00", X"75", X"53", X"00", X"71", X"0a", 
    X"80", X"14", X"e5", X"81", X"b4", X"51", X"0f", X"e5", 
    X"50", X"b4", X"08", X"0a", X"e5", X"51", X"b4", X"23", 
    X"05", X"75", X"99", X"61", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"12", X"80", X"0c", X"80", 
    X"06", X"00", X"75", X"99", X"62", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"90", X"7f", X"cd", 
    X"74", X"33", X"73", X"02", X"23", X"4d", X"00", X"00", 
    X"74", X"00", X"74", X"00", X"74", X"00", X"74", X"00", 
    X"75", X"99", X"63", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"02", X"80", X"06", X"02", X"23", 
    X"62", X"00", X"00", X"00", X"00", X"75", X"99", X"64", 
    X"80", X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", 
    X"74", X"00", X"61", X"6e", X"80", X"02", X"74", X"42", 
    X"b4", X"42", X"06", X"00", X"75", X"99", X"65", X"80", 
    X"06", X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", 
    X"99", X"0d", X"75", X"99", X"0a", X"75", X"99", X"53", 
    X"75", X"81", X"4f", X"75", X"4f", X"23", X"75", X"4e", 
    X"9c", X"75", X"4d", X"23", X"75", X"4c", X"a6", X"22", 
    X"80", X"16", X"74", X"00", X"e5", X"81", X"b4", X"4d", 
    X"0f", X"22", X"80", X"0c", X"74", X"00", X"e5", X"81", 
    X"b4", X"4b", X"05", X"75", X"99", X"61", X"80", X"06", 
    X"75", X"99", X"3f", X"75", X"6e", X"01", X"75", X"81", 
    X"4f", X"75", X"4f", X"23", X"75", X"4e", X"ca", X"75", 
    X"4d", X"23", X"75", X"4c", X"d4", X"22", X"80", X"e8", 
    X"74", X"00", X"e5", X"81", X"b4", X"4d", X"0f", X"22", 
    X"80", X"de", X"74", X"00", X"e5", X"81", X"b4", X"4b", 
    X"05", X"75", X"99", X"62", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"75", X"99", X"0d", X"75", 
    X"99", X"0a", X"75", X"99", X"54", X"75", X"f0", X"07", 
    X"74", X"13", X"e5", X"f0", X"b4", X"07", X"37", X"90", 
    X"24", X"36", X"78", X"00", X"79", X"09", X"e8", X"08", 
    X"93", X"f5", X"f0", X"e8", X"08", X"93", X"84", X"f5", 
    X"60", X"e8", X"08", X"93", X"70", X"15", X"e5", X"d0", 
    X"54", X"04", X"70", X"1a", X"e8", X"08", X"93", X"b5", 
    X"60", X"14", X"e8", X"08", X"93", X"b5", X"f0", X"0e", 
    X"02", X"24", X"25", X"08", X"08", X"19", X"e9", X"70", 
    X"d5", X"75", X"99", X"61", X"80", X"06", X"75", X"99", 
    X"3f", X"75", X"6e", X"01", X"80", X"2d", X"07", X"13", 
    X"00", X"02", X"05", X"07", X"11", X"00", X"02", X"03", 
    X"07", X"0d", X"00", X"01", X"06", X"0d", X"11", X"00", 
    X"01", X"04", X"11", X"0d", X"00", X"00", X"0d", X"00", 
    X"0d", X"04", X"00", X"0d", X"80", X"87", X"00", X"01", 
    X"07", X"01", X"ff", X"00", X"ff", X"00", X"02", X"ff", 
    X"00", X"7f", X"01", X"90", X"24", X"a4", X"78", X"00", 
    X"79", X"09", X"e8", X"08", X"93", X"f5", X"f0", X"e8", 
    X"08", X"93", X"a4", X"f5", X"60", X"e8", X"93", X"60", 
    X"08", X"e5", X"d0", X"54", X"04", X"60", X"1d", X"80", 
    X"06", X"e5", X"d0", X"54", X"04", X"70", X"15", X"e8", 
    X"08", X"93", X"b5", X"f0", X"0f", X"e8", X"08", X"93", 
    X"b5", X"60", X"09", X"19", X"e9", X"70", X"d3", X"75", 
    X"99", X"62", X"80", X"06", X"75", X"99", X"3f", X"75", 
    X"6e", X"01", X"80", X"24", X"07", X"13", X"00", X"85", 
    X"07", X"11", X"00", X"77", X"07", X"0d", X"00", X"5b", 
    X"0d", X"11", X"00", X"dd", X"11", X"0d", X"00", X"dd", 
    X"00", X"0d", X"00", X"00", X"80", X"87", X"43", X"80", 
    X"01", X"ff", X"00", X"ff", X"02", X"ff", X"01", X"fe", 
    X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", X"99", 
    X"55", X"75", X"d0", X"00", X"74", X"01", X"12", X"24", 
    X"f3", X"75", X"d0", X"08", X"74", X"09", X"12", X"24", 
    X"f3", X"75", X"d0", X"10", X"74", X"11", X"12", X"24", 
    X"f3", X"75", X"d0", X"18", X"74", X"19", X"12", X"24", 
    X"f3", X"80", X"1e", X"f8", X"79", X"12", X"7f", X"34", 
    X"e6", X"b4", X"12", X"1b", X"74", X"56", X"f6", X"b9", 
    X"56", X"15", X"e8", X"24", X"06", X"f8", X"e6", X"b4", 
    X"34", X"0d", X"74", X"78", X"f6", X"b4", X"78", X"07", 
    X"22", X"00", X"75", X"99", X"61", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", X"0d", 
    X"75", X"99", X"0a", X"75", X"99", X"56", X"a5", X"00", 
    X"75", X"99", X"61", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"75", X"d0", X"00", X"74", X"1a", 
    X"d4", X"85", X"d0", X"70", X"b4", X"20", X"4e", X"e5", 
    X"70", X"b4", X"01", X"49", X"75", X"d0", X"40", X"74", 
    X"12", X"d4", X"85", X"d0", X"70", X"b4", X"18", X"3d", 
    X"e5", X"70", X"b4", X"40", X"38", X"75", X"d0", X"40", 
    X"74", X"1a", X"d4", X"85", X"d0", X"70", X"b4", X"20", 
    X"2c", X"e5", X"70", X"b4", X"41", X"27", X"75", X"d0", 
    X"c0", X"74", X"00", X"d4", X"85", X"d0", X"70", X"b4", 
    X"66", X"1b", X"e5", X"70", X"b4", X"c0", X"16", X"75", 
    X"d0", X"40", X"74", X"fa", X"d4", X"85", X"d0", X"70", 
    X"b4", X"60", X"0a", X"e5", X"70", X"b4", X"c0", X"05", 
    X"75", X"99", X"62", X"80", X"06", X"75", X"99", X"3f", 
    X"75", X"6e", X"01", X"78", X"31", X"79", X"32", X"74", 
    X"42", X"f6", X"04", X"f7", X"74", X"76", X"d6", X"b4", 
    X"72", X"15", X"e5", X"31", X"b4", X"46", X"10", X"74", 
    X"79", X"d7", X"b4", X"73", X"0a", X"e5", X"32", X"b4", 
    X"49", X"05", X"75", X"99", X"63", X"80", X"06", X"75", 
    X"99", X"3f", X"75", X"6e", X"01", X"75", X"99", X"0d", 
    X"75", X"99", X"0a", X"e5", X"6e", X"70", X"1a", X"75", 
    X"99", X"0d", X"75", X"99", X"0a", X"75", X"99", X"50", 
    X"75", X"99", X"41", X"75", X"99", X"53", X"75", X"99", 
    X"53", X"75", X"99", X"0d", X"75", X"99", X"0a", X"80", 
    X"1a", X"75", X"99", X"0d", X"75", X"99", X"0a", X"75", 
    X"99", X"46", X"75", X"99", X"41", X"75", X"99", X"49", 
    X"75", X"99", X"4c", X"75", X"99", X"0d", X"75", X"99", 
    X"0a", X"80", X"00", X"75", X"99", X"04", X"a1", X"fe", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"02", X"23", X"40", X"02", X"23", X"4d", X"02", X"23", 
    X"5b", X"02", X"23", X"62", X"e5", X"81", X"b4", X"53", 
    X"0d", X"e5", X"52", X"b4", X"27", X"08", X"e5", X"53", 
    X"b4", X"23", X"03", X"02", X"23", X"29", X"02", X"23", 
    X"2f" 
);


end package obj_code_pkg;
