--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- This is where the application code lives.
-- FIXME should only be used from top level entity
-- FIXME name of package should be application-related
-- FIXME convert to vhdl template
--------------------------------------------------------------------------------
-- Copyright (C) 2011 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.light52_pkg.all;

package obj_code_pkg is

constant object_code : t_obj_code(0 to 10107) := (
    X"02", X"00", X"13", X"32", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"02", X"15", X"4e", X"12", X"00", 
    X"81", X"80", X"fe", X"75", X"81", X"3a", X"12", X"22", 
    X"6b", X"e5", X"82", X"60", X"03", X"02", X"00", X"0e", 
    X"79", X"1a", X"e9", X"44", X"00", X"60", X"1b", X"7a", 
    X"01", X"90", X"27", X"62", X"78", X"8c", X"75", X"a0", 
    X"06", X"e4", X"93", X"f2", X"a3", X"08", X"b8", X"00", 
    X"02", X"05", X"a0", X"d9", X"f4", X"da", X"f2", X"75", 
    X"a0", X"ff", X"e4", X"78", X"ff", X"f6", X"d8", X"fd", 
    X"78", X"00", X"e8", X"44", X"00", X"60", X"0a", X"79", 
    X"00", X"75", X"a0", X"00", X"e4", X"f3", X"09", X"d8", 
    X"fc", X"78", X"8c", X"e8", X"44", X"06", X"60", X"0c", 
    X"79", X"07", X"90", X"00", X"00", X"e4", X"f0", X"a3", 
    X"d8", X"fc", X"d9", X"fa", X"90", X"06", X"1a", X"74", 
    X"b6", X"f0", X"a3", X"74", X"05", X"f0", X"a3", X"e4", 
    X"f0", X"90", X"06", X"2f", X"e4", X"f0", X"02", X"00", 
    X"0e", X"12", X"14", X"21", X"90", X"06", X"20", X"74", 
    X"78", X"f0", X"a3", X"74", X"22", X"f0", X"a3", X"74", 
    X"80", X"f0", X"90", X"22", X"6f", X"75", X"f0", X"80", 
    X"12", X"13", X"e8", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"ed", X"4e", X"70", X"1b", X"74", X"7b", X"c0", 
    X"e0", X"74", X"22", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"90", X"00", X"01", X"12", X"13", X"e4", 
    X"90", X"00", X"26", X"12", X"13", X"86", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"90", X"00", X"03", X"ed", 
    X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"90", 
    X"00", X"26", X"12", X"13", X"86", X"ad", X"82", X"ae", 
    X"83", X"af", X"f0", X"90", X"00", X"00", X"ed", X"f0", 
    X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"90", X"00", 
    X"03", X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", 
    X"fc", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"ea", 
    X"12", X"17", X"7d", X"a3", X"eb", X"12", X"17", X"7d", 
    X"a3", X"ec", X"12", X"17", X"7d", X"74", X"03", X"2d", 
    X"fa", X"e4", X"3e", X"fb", X"8f", X"04", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"e4", X"12", X"17", X"7d", 
    X"74", X"04", X"2d", X"fa", X"e4", X"3e", X"fb", X"8f", 
    X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"74", 
    X"02", X"12", X"17", X"7d", X"74", X"05", X"2d", X"fa", 
    X"e4", X"3e", X"fb", X"8f", X"04", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"74", X"28", X"12", X"17", X"7d", 
    X"a3", X"e4", X"12", X"17", X"7d", X"74", X"07", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"90", X"06", X"31", X"74", 
    X"93", X"f0", X"a3", X"74", X"22", X"f0", X"a3", X"74", 
    X"80", X"f0", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"15", X"a5", X"90", X"06", X"31", X"74", X"b2", 
    X"f0", X"a3", X"74", X"22", X"f0", X"a3", X"74", X"80", 
    X"f0", X"90", X"05", X"4b", X"75", X"f0", X"00", X"12", 
    X"15", X"a5", X"90", X"01", X"dc", X"74", X"0a", X"f0", 
    X"a3", X"e4", X"f0", X"74", X"d1", X"c0", X"e0", X"74", 
    X"22", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"1a", X"0b", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"74", X"d3", X"c0", X"e0", X"74", X"22", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"74", X"d1", X"c0", 
    X"e0", X"74", X"22", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"74", X"a8", X"c0", X"e0", X"74", X"61", 
    X"c0", X"e0", X"74", X"03", X"c0", X"e0", X"74", X"23", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", X"12", 
    X"14", X"44", X"ac", X"82", X"ad", X"83", X"ae", X"f0", 
    X"ff", X"90", X"05", X"20", X"ec", X"f0", X"a3", X"ed", 
    X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"7e", 
    X"01", X"7f", X"00", X"c3", X"74", X"a8", X"9e", X"74", 
    X"e1", X"8f", X"f0", X"63", X"f0", X"80", X"95", X"f0", 
    X"50", X"03", X"02", X"04", X"81", X"c0", X"07", X"c0", 
    X"06", X"12", X"0f", X"63", X"12", X"0f", X"3b", X"90", 
    X"05", X"44", X"74", X"02", X"f0", X"a3", X"e4", X"f0", 
    X"90", X"05", X"46", X"74", X"03", X"f0", X"a3", X"e4", 
    X"f0", X"90", X"06", X"31", X"74", X"30", X"f0", X"a3", 
    X"74", X"23", X"f0", X"a3", X"74", X"80", X"f0", X"90", 
    X"05", X"6a", X"75", X"f0", X"00", X"12", X"15", X"a5", 
    X"90", X"05", X"4a", X"74", X"01", X"f0", X"90", X"05", 
    X"aa", X"74", X"6a", X"f0", X"a3", X"74", X"05", X"f0", 
    X"a3", X"e4", X"f0", X"90", X"05", X"4b", X"75", X"f0", 
    X"00", X"12", X"12", X"4d", X"ac", X"82", X"ad", X"83", 
    X"d0", X"06", X"d0", X"07", X"ec", X"4d", X"b4", X"01", 
    X"00", X"e4", X"33", X"fc", X"90", X"00", X"08", X"f0", 
    X"ec", X"33", X"95", X"e0", X"a3", X"f0", X"7c", X"02", 
    X"7d", X"00", X"c3", X"ec", X"94", X"03", X"ed", X"64", 
    X"80", X"94", X"80", X"50", X"67", X"90", X"06", X"4c", 
    X"ec", X"f0", X"a3", X"ed", X"f0", X"90", X"00", X"05", 
    X"c0", X"07", X"c0", X"06", X"c0", X"05", X"c0", X"04", 
    X"12", X"17", X"96", X"e5", X"82", X"85", X"83", X"f0", 
    X"d0", X"04", X"d0", X"05", X"24", X"fd", X"fa", X"e5", 
    X"f0", X"34", X"ff", X"fb", X"90", X"05", X"48", X"ea", 
    X"f0", X"a3", X"eb", X"f0", X"90", X"05", X"97", X"74", 
    X"03", X"f0", X"a3", X"e4", X"f0", X"90", X"05", X"99", 
    X"74", X"48", X"f0", X"a3", X"74", X"05", X"f0", X"a3", 
    X"e4", X"f0", X"8c", X"82", X"8d", X"83", X"c0", X"05", 
    X"c0", X"04", X"12", X"10", X"24", X"d0", X"04", X"d0", 
    X"05", X"d0", X"06", X"d0", X"07", X"0c", X"bc", X"00", 
    X"01", X"0d", X"90", X"05", X"44", X"ec", X"f0", X"a3", 
    X"ed", X"f0", X"80", X"8e", X"90", X"05", X"44", X"ec", 
    X"f0", X"a3", X"ed", X"f0", X"90", X"05", X"48", X"e0", 
    X"fa", X"a3", X"e0", X"fb", X"90", X"05", X"9e", X"74", 
    X"3e", X"f0", X"a3", X"74", X"00", X"f0", X"a3", X"e4", 
    X"f0", X"90", X"05", X"a1", X"ec", X"f0", X"a3", X"ed", 
    X"f0", X"90", X"05", X"a3", X"ea", X"f0", X"a3", X"eb", 
    X"f0", X"90", X"00", X"0c", X"75", X"f0", X"00", X"c0", 
    X"07", X"c0", X"06", X"12", X"10", X"66", X"90", X"00", 
    X"00", X"e0", X"fb", X"a3", X"e0", X"fc", X"a3", X"e0", 
    X"fd", X"8b", X"82", X"8c", X"83", X"8d", X"f0", X"12", 
    X"0c", X"2b", X"d0", X"06", X"d0", X"07", X"8e", X"04", 
    X"8f", X"05", X"7b", X"41", X"90", X"00", X"0b", X"e0", 
    X"fa", X"c3", X"64", X"80", X"8b", X"f0", X"63", X"f0", 
    X"80", X"95", X"f0", X"40", X"7b", X"90", X"05", X"a8", 
    X"74", X"43", X"f0", X"8b", X"82", X"c0", X"07", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", X"12", 
    X"12", X"2e", X"aa", X"82", X"d0", X"03", X"d0", X"04", 
    X"d0", X"05", X"d0", X"06", X"d0", X"07", X"90", X"05", 
    X"4a", X"e0", X"f9", X"b5", X"02", X"4e", X"90", X"05", 
    X"93", X"74", X"4a", X"f0", X"a3", X"74", X"05", X"f0", 
    X"a3", X"e4", X"f0", X"75", X"82", X"00", X"c0", X"07", 
    X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", 
    X"12", X"0f", X"71", X"90", X"06", X"31", X"74", X"4f", 
    X"f0", X"a3", X"74", X"23", X"f0", X"a3", X"74", X"80", 
    X"f0", X"90", X"05", X"6a", X"75", X"f0", X"00", X"12", 
    X"15", X"a5", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"d0", X"07", X"90", X"05", X"46", X"ec", 
    X"f0", X"a3", X"ed", X"f0", X"90", X"00", X"06", X"ec", 
    X"f0", X"a3", X"ed", X"f0", X"0b", X"02", X"03", X"4c", 
    X"90", X"05", X"44", X"e0", X"fc", X"a3", X"e0", X"fd", 
    X"90", X"05", X"46", X"e0", X"fa", X"a3", X"e0", X"fb", 
    X"90", X"06", X"4c", X"ec", X"f0", X"a3", X"ed", X"f0", 
    X"8a", X"82", X"8b", X"83", X"c0", X"07", X"c0", X"06", 
    X"12", X"17", X"96", X"e5", X"82", X"85", X"83", X"f0", 
    X"90", X"05", X"46", X"f0", X"a3", X"e5", X"f0", X"f0", 
    X"90", X"05", X"48", X"e0", X"fc", X"a3", X"e0", X"fd", 
    X"90", X"05", X"46", X"e0", X"fa", X"a3", X"e0", X"fb", 
    X"90", X"06", X"58", X"ec", X"f0", X"a3", X"ed", X"f0", 
    X"8a", X"82", X"8b", X"83", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"c0", X"02", X"12", X"18", X"b6", X"a8", 
    X"82", X"a9", X"83", X"d0", X"02", X"d0", X"03", X"d0", 
    X"04", X"d0", X"05", X"90", X"05", X"44", X"e8", X"f0", 
    X"a3", X"e9", X"f0", X"90", X"06", X"4c", X"ea", X"c3", 
    X"9c", X"f0", X"eb", X"9d", X"a3", X"f0", X"90", X"00", 
    X"07", X"c0", X"01", X"c0", X"00", X"12", X"17", X"96", 
    X"e5", X"82", X"85", X"83", X"f0", X"d0", X"00", X"d0", 
    X"01", X"90", X"05", X"46", X"c3", X"98", X"f0", X"e5", 
    X"f0", X"99", X"a3", X"f0", X"90", X"05", X"44", X"75", 
    X"f0", X"00", X"12", X"0e", X"4d", X"d0", X"06", X"d0", 
    X"07", X"0e", X"be", X"00", X"01", X"0f", X"02", X"02", 
    X"03", X"12", X"14", X"44", X"ac", X"82", X"ad", X"83", 
    X"ae", X"f0", X"ff", X"90", X"05", X"24", X"ec", X"f0", 
    X"a3", X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", 
    X"f0", X"74", X"6e", X"c0", X"e0", X"74", X"23", X"c0", 
    X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"74", X"d1", 
    X"c0", X"e0", X"74", X"22", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"74", X"7e", X"c0", X"e0", X"74", 
    X"23", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"1a", X"0b", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"74", X"d1", X"c0", X"e0", X"74", X"22", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"90", X"00", X"06", 
    X"e0", X"c0", X"e0", X"a3", X"e0", X"c0", X"e0", X"74", 
    X"b4", X"c0", X"e0", X"74", X"23", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", 
    X"24", X"fb", X"f5", X"81", X"74", X"05", X"c0", X"e0", 
    X"e4", X"c0", X"e0", X"74", X"cd", X"c0", X"e0", X"74", 
    X"23", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", 
    X"90", X"00", X"08", X"e0", X"c0", X"e0", X"a3", X"e0", 
    X"c0", X"e0", X"74", X"e6", X"c0", X"e0", X"74", X"23", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", X"74", 
    X"01", X"c0", X"e0", X"e4", X"c0", X"e0", X"74", X"cd", 
    X"c0", X"e0", X"74", X"23", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"90", X"00", X"0a", X"e0", X"ff", 
    X"33", X"95", X"e0", X"fe", X"c0", X"07", X"c0", X"06", 
    X"74", X"ff", X"c0", X"e0", X"74", X"23", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", 
    X"81", X"24", X"fb", X"f5", X"81", X"74", X"41", X"c0", 
    X"e0", X"e4", X"c0", X"e0", X"74", X"18", X"c0", X"e0", 
    X"74", X"24", X"c0", X"e0", X"74", X"80", X"c0", X"e0", 
    X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", 
    X"81", X"90", X"00", X"0b", X"e0", X"ff", X"33", X"95", 
    X"e0", X"fe", X"c0", X"07", X"c0", X"06", X"74", X"31", 
    X"c0", X"e0", X"74", X"24", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"74", X"42", X"c0", X"e0", X"e4", 
    X"c0", X"e0", X"74", X"18", X"c0", X"e0", X"74", X"24", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", X"90", 
    X"00", X"1c", X"e0", X"fe", X"a3", X"e0", X"ff", X"c0", 
    X"06", X"c0", X"07", X"74", X"4a", X"c0", X"e0", X"74", 
    X"24", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", 
    X"74", X"07", X"c0", X"e0", X"e4", X"c0", X"e0", X"74", 
    X"cd", X"c0", X"e0", X"74", X"23", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", 
    X"24", X"fb", X"f5", X"81", X"90", X"01", X"dc", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"c0", X"06", X"c0", X"07", 
    X"74", X"63", X"c0", X"e0", X"74", X"24", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", 
    X"81", X"24", X"fb", X"f5", X"81", X"74", X"7c", X"c0", 
    X"e0", X"74", X"24", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"74", X"a6", X"c0", X"e0", X"74", X"24", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"15", X"81", X"15", X"81", X"15", X"81", X"90", 
    X"00", X"00", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"22", X"4f", X"fd", X"a3", X"12", X"22", X"4f", 
    X"fe", X"a3", X"12", X"22", X"4f", X"c0", X"05", X"c0", 
    X"06", X"74", X"b2", X"c0", X"e0", X"74", X"24", X"c0", 
    X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", 
    X"e5", X"81", X"24", X"fb", X"f5", X"81", X"74", X"cb", 
    X"c0", X"e0", X"74", X"24", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"90", X"00", X"00", X"e0", X"fd", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"03", 
    X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"22", X"4f", X"fd", X"7f", 
    X"00", X"c0", X"05", X"c0", X"07", X"74", X"fc", X"c0", 
    X"e0", X"74", X"24", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", 
    X"f5", X"81", X"e4", X"c0", X"e0", X"c0", X"e0", X"74", 
    X"cd", X"c0", X"e0", X"74", X"23", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", 
    X"24", X"fb", X"f5", X"81", X"90", X"00", X"00", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", 
    X"04", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"22", X"4f", X"fd", 
    X"7f", X"00", X"c0", X"05", X"c0", X"07", X"74", X"15", 
    X"c0", X"e0", X"74", X"25", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"74", X"02", X"c0", X"e0", X"e4", 
    X"c0", X"e0", X"74", X"cd", X"c0", X"e0", X"74", X"23", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", X"90", 
    X"00", X"00", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"74", X"05", X"2d", X"fd", X"e4", X"3e", 
    X"fe", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"22", X"4f", X"fd", X"a3", X"12", X"22", X"4f", X"fe", 
    X"c0", X"05", X"c0", X"06", X"74", X"2e", X"c0", X"e0", 
    X"74", X"25", X"c0", X"e0", X"74", X"80", X"c0", X"e0", 
    X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", 
    X"81", X"74", X"11", X"c0", X"e0", X"e4", X"c0", X"e0", 
    X"74", X"cd", X"c0", X"e0", X"74", X"23", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", 
    X"81", X"24", X"fb", X"f5", X"81", X"90", X"00", X"00", 
    X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"74", X"07", X"2d", X"fd", X"e4", X"3e", X"fe", X"c0", 
    X"05", X"c0", X"06", X"c0", X"07", X"74", X"47", X"c0", 
    X"e0", X"74", X"25", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fa", 
    X"f5", X"81", X"74", X"60", X"c0", X"e0", X"74", X"25", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"15", X"81", X"15", X"81", X"15", X"81", X"74", 
    X"95", X"c0", X"e0", X"74", X"25", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"15", X"81", 
    X"15", X"81", X"15", X"81", X"90", X"00", X"03", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"22", X"4f", 
    X"fd", X"a3", X"12", X"22", X"4f", X"fe", X"a3", X"12", 
    X"22", X"4f", X"c0", X"05", X"c0", X"06", X"74", X"b2", 
    X"c0", X"e0", X"74", X"24", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"74", X"a6", X"c0", X"e0", X"74", 
    X"25", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"1a", X"0b", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"90", X"00", X"03", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"74", X"03", X"2d", X"fd", X"e4", 
    X"3e", X"fe", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"22", X"4f", X"fd", X"7f", X"00", X"c0", X"05", 
    X"c0", X"07", X"74", X"fc", X"c0", X"e0", X"74", X"24", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", X"e4", 
    X"c0", X"e0", X"c0", X"e0", X"74", X"cd", X"c0", X"e0", 
    X"74", X"23", X"c0", X"e0", X"74", X"80", X"c0", X"e0", 
    X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", 
    X"81", X"90", X"00", X"03", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"74", X"04", X"2d", X"fd", 
    X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"22", X"4f", X"fd", X"7f", X"00", X"c0", 
    X"05", X"c0", X"07", X"74", X"15", X"c0", X"e0", X"74", 
    X"25", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", 
    X"74", X"01", X"c0", X"e0", X"e4", X"c0", X"e0", X"74", 
    X"cd", X"c0", X"e0", X"74", X"23", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", 
    X"24", X"fb", X"f5", X"81", X"90", X"00", X"03", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", 
    X"05", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"22", X"4f", X"fd", 
    X"a3", X"12", X"22", X"4f", X"fe", X"c0", X"05", X"c0", 
    X"06", X"74", X"2e", X"c0", X"e0", X"74", X"25", X"c0", 
    X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", 
    X"e5", X"81", X"24", X"fb", X"f5", X"81", X"74", X"12", 
    X"c0", X"e0", X"e4", X"c0", X"e0", X"74", X"cd", X"c0", 
    X"e0", X"74", X"23", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", 
    X"f5", X"81", X"90", X"00", X"03", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"07", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"74", X"47", X"c0", X"e0", X"74", X"25", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"e5", X"81", X"24", X"fa", X"f5", X"81", X"74", 
    X"60", X"c0", X"e0", X"74", X"25", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"15", X"81", 
    X"15", X"81", X"15", X"81", X"90", X"05", X"44", X"e0", 
    X"c0", X"e0", X"a3", X"e0", X"c0", X"e0", X"74", X"e6", 
    X"c0", X"e0", X"74", X"25", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"74", X"05", X"c0", X"e0", X"e4", 
    X"c0", X"e0", X"74", X"cd", X"c0", X"e0", X"74", X"23", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"e5", X"81", X"24", X"fb", X"f5", X"81", X"90", 
    X"05", X"46", X"e0", X"c0", X"e0", X"a3", X"e0", X"c0", 
    X"e0", X"74", X"ff", X"c0", X"e0", X"74", X"25", X"c0", 
    X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", 
    X"e5", X"81", X"24", X"fb", X"f5", X"81", X"74", X"0d", 
    X"c0", X"e0", X"e4", X"c0", X"e0", X"74", X"cd", X"c0", 
    X"e0", X"74", X"23", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", 
    X"f5", X"81", X"90", X"05", X"48", X"e0", X"c0", X"e0", 
    X"a3", X"e0", X"c0", X"e0", X"74", X"18", X"c0", X"e0", 
    X"74", X"26", X"c0", X"e0", X"74", X"80", X"c0", X"e0", 
    X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", 
    X"81", X"74", X"07", X"c0", X"e0", X"e4", X"c0", X"e0", 
    X"74", X"cd", X"c0", X"e0", X"74", X"23", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", 
    X"81", X"24", X"fb", X"f5", X"81", X"90", X"05", X"4a", 
    X"e0", X"ff", X"7e", X"00", X"c0", X"07", X"c0", X"06", 
    X"74", X"31", X"c0", X"e0", X"74", X"26", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", 
    X"81", X"24", X"fb", X"f5", X"81", X"74", X"01", X"c0", 
    X"e0", X"e4", X"c0", X"e0", X"74", X"cd", X"c0", X"e0", 
    X"74", X"23", X"c0", X"e0", X"74", X"80", X"c0", X"e0", 
    X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", X"f5", 
    X"81", X"74", X"4b", X"c0", X"e0", X"74", X"05", X"c0", 
    X"e0", X"e4", X"c0", X"e0", X"74", X"4a", X"c0", X"e0", 
    X"74", X"26", X"c0", X"e0", X"74", X"80", X"c0", X"e0", 
    X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fa", X"f5", 
    X"81", X"74", X"63", X"c0", X"e0", X"74", X"26", X"c0", 
    X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"74", X"6a", 
    X"c0", X"e0", X"74", X"05", X"c0", X"e0", X"e4", X"c0", 
    X"e0", X"74", X"98", X"c0", X"e0", X"74", X"26", X"c0", 
    X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", 
    X"e5", X"81", X"24", X"fa", X"f5", X"81", X"74", X"b1", 
    X"c0", X"e0", X"74", X"26", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"1a", X"0b", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"74", X"d1", X"c0", X"e0", X"74", 
    X"22", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"1a", X"0b", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"90", X"05", X"20", X"e0", X"fc", X"a3", X"e0", X"fd", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"90", X"05", 
    X"24", X"e0", X"f8", X"a3", X"e0", X"f9", X"a3", X"e0", 
    X"fa", X"a3", X"e0", X"fb", X"90", X"05", X"24", X"e8", 
    X"c3", X"9c", X"f0", X"e9", X"9d", X"a3", X"f0", X"ea", 
    X"9e", X"a3", X"f0", X"eb", X"9f", X"a3", X"f0", X"90", 
    X"05", X"24", X"e0", X"fc", X"a3", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"90", X"06", X"37", 
    X"74", X"e8", X"f0", X"a3", X"74", X"03", X"f0", X"a3", 
    X"e4", X"f0", X"a3", X"f0", X"8c", X"82", X"8d", X"83", 
    X"8e", X"f0", X"ef", X"c0", X"07", X"c0", X"06", X"c0", 
    X"05", X"c0", X"04", X"12", X"15", X"fe", X"85", X"82", 
    X"08", X"85", X"83", X"09", X"85", X"f0", X"0a", X"f5", 
    X"0b", X"90", X"06", X"54", X"e5", X"08", X"f0", X"a3", 
    X"e5", X"09", X"f0", X"a3", X"e5", X"0a", X"f0", X"a3", 
    X"e5", X"0b", X"f0", X"90", X"03", X"e8", X"e4", X"f5", 
    X"f0", X"12", X"18", X"4a", X"a8", X"82", X"a9", X"83", 
    X"aa", X"f0", X"fb", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"d0", X"07", X"ec", X"c3", X"98", X"fc", X"ed", 
    X"99", X"fd", X"ee", X"9a", X"fe", X"ef", X"9b", X"ff", 
    X"c0", X"04", X"c0", X"05", X"c0", X"06", X"c0", X"07", 
    X"c0", X"08", X"c0", X"09", X"c0", X"0a", X"c0", X"0b", 
    X"74", X"e6", X"c0", X"e0", X"74", X"26", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"1a", X"0b", X"e5", 
    X"81", X"24", X"f5", X"f5", X"81", X"90", X"05", X"24", 
    X"e0", X"fc", X"a3", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"90", X"06", X"37", X"ec", X"f0", 
    X"a3", X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", 
    X"f0", X"90", X"78", X"40", X"75", X"f0", X"7d", X"74", 
    X"01", X"12", X"15", X"fe", X"ac", X"82", X"ad", X"83", 
    X"ae", X"f0", X"ff", X"90", X"05", X"28", X"ec", X"f0", 
    X"a3", X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", 
    X"f0", X"c0", X"04", X"c0", X"05", X"74", X"10", X"c0", 
    X"e0", X"74", X"27", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"1a", X"0b", X"e5", X"81", X"24", X"fb", 
    X"f5", X"81", X"74", X"2c", X"c0", X"e0", X"74", X"27", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"1a", 
    X"0b", X"15", X"81", X"15", X"81", X"15", X"81", X"90", 
    X"00", X"00", X"22", X"af", X"f0", X"ae", X"83", X"e5", 
    X"82", X"90", X"05", X"89", X"f0", X"a3", X"ee", X"f0", 
    X"a3", X"ef", X"f0", X"90", X"05", X"89", X"e0", X"f5", 
    X"0c", X"a3", X"e0", X"f5", X"0d", X"a3", X"e0", X"f5", 
    X"0e", X"85", X"0c", X"82", X"85", X"0d", X"83", X"85", 
    X"0e", X"f0", X"12", X"22", X"4f", X"fa", X"a3", X"12", 
    X"22", X"4f", X"fb", X"a3", X"12", X"22", X"4f", X"fc", 
    X"8a", X"00", X"8b", X"01", X"8c", X"07", X"88", X"0f", 
    X"89", X"10", X"8f", X"11", X"90", X"00", X"00", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"90", 
    X"06", X"43", X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", 
    X"ef", X"f0", X"90", X"06", X"46", X"74", X"26", X"f0", 
    X"a3", X"e4", X"f0", X"85", X"0f", X"82", X"85", X"10", 
    X"83", X"85", X"11", X"f0", X"c0", X"04", X"c0", X"03", 
    X"c0", X"02", X"12", X"17", X"09", X"d0", X"02", X"d0", 
    X"03", X"d0", X"04", X"74", X"04", X"25", X"0c", X"f5", 
    X"0f", X"e4", X"35", X"0d", X"f5", X"10", X"85", X"0e", 
    X"11", X"74", X"05", X"25", X"0c", X"f5", X"12", X"e4", 
    X"35", X"0d", X"f5", X"13", X"85", X"0e", X"14", X"85", 
    X"12", X"82", X"85", X"13", X"83", X"85", X"14", X"f0", 
    X"74", X"05", X"12", X"17", X"7d", X"a3", X"e4", X"12", 
    X"17", X"7d", X"74", X"04", X"2a", X"fd", X"e4", X"3b", 
    X"fe", X"8c", X"07", X"0d", X"bd", X"00", X"01", X"0e", 
    X"85", X"12", X"82", X"85", X"13", X"83", X"85", X"14", 
    X"f0", X"12", X"22", X"4f", X"f8", X"a3", X"12", X"22", 
    X"4f", X"f9", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e8", X"12", X"17", X"7d", X"a3", X"e9", X"12", X"17", 
    X"7d", X"85", X"0c", X"82", X"85", X"0d", X"83", X"85", 
    X"0e", X"f0", X"12", X"22", X"4f", X"fd", X"a3", X"12", 
    X"22", X"4f", X"fe", X"a3", X"12", X"22", X"4f", X"ff", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"ed", X"12", 
    X"17", X"7d", X"a3", X"ee", X"12", X"17", X"7d", X"a3", 
    X"ef", X"12", X"17", X"7d", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"c0", X"04", X"c0", X"03", X"c0", X"02", 
    X"12", X"0e", X"b6", X"d0", X"02", X"d0", X"03", X"d0", 
    X"04", X"74", X"03", X"2a", X"fd", X"e4", X"3b", X"fe", 
    X"8c", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"22", X"4f", X"60", X"03", X"02", X"0e", X"13", 
    X"74", X"04", X"2a", X"f5", X"12", X"e4", X"3b", X"f5", 
    X"13", X"8c", X"14", X"74", X"01", X"25", X"12", X"f8", 
    X"e4", X"35", X"13", X"f9", X"af", X"14", X"88", X"82", 
    X"89", X"83", X"8f", X"f0", X"74", X"06", X"12", X"17", 
    X"7d", X"a3", X"e4", X"12", X"17", X"7d", X"85", X"0f", 
    X"82", X"85", X"10", X"83", X"85", X"11", X"f0", X"12", 
    X"22", X"4f", X"ff", X"90", X"05", X"93", X"e5", X"12", 
    X"f0", X"a3", X"e5", X"13", X"f0", X"a3", X"e5", X"14", 
    X"f0", X"8f", X"82", X"c0", X"04", X"c0", X"03", X"c0", 
    X"02", X"12", X"0f", X"71", X"d0", X"02", X"d0", X"03", 
    X"d0", X"04", X"90", X"00", X"00", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"22", X"4f", X"fd", X"a3", 
    X"12", X"22", X"4f", X"fe", X"a3", X"12", X"22", X"4f", 
    X"ff", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"ed", 
    X"12", X"17", X"7d", X"a3", X"ee", X"12", X"17", X"7d", 
    X"a3", X"ef", X"12", X"17", X"7d", X"74", X"04", X"2a", 
    X"fa", X"e4", X"3b", X"fb", X"0a", X"ba", X"00", X"01", 
    X"0b", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", 
    X"22", X"4f", X"fe", X"a3", X"12", X"22", X"4f", X"ff", 
    X"90", X"05", X"97", X"74", X"0a", X"f0", X"a3", X"e4", 
    X"f0", X"90", X"05", X"99", X"ea", X"f0", X"a3", X"eb", 
    X"f0", X"a3", X"ec", X"f0", X"8e", X"82", X"8f", X"83", 
    X"02", X"10", X"24", X"ad", X"0c", X"ae", X"0d", X"af", 
    X"0e", X"85", X"0c", X"82", X"85", X"0d", X"83", X"85", 
    X"0e", X"f0", X"12", X"22", X"4f", X"fa", X"a3", X"12", 
    X"22", X"4f", X"fb", X"a3", X"12", X"22", X"4f", X"fc", 
    X"90", X"06", X"43", X"ea", X"f0", X"a3", X"eb", X"f0", 
    X"a3", X"ec", X"f0", X"90", X"06", X"46", X"74", X"26", 
    X"f0", X"a3", X"e4", X"f0", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"02", X"17", X"09", X"af", X"f0", X"ae", 
    X"83", X"e5", X"82", X"90", X"05", X"8c", X"f0", X"a3", 
    X"ee", X"f0", X"a3", X"ef", X"f0", X"90", X"05", X"8c", 
    X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"22", 
    X"4f", X"fb", X"a3", X"12", X"22", X"4f", X"fc", X"74", 
    X"0a", X"2b", X"fb", X"e4", X"3c", X"fc", X"90", X"00", 
    X"0a", X"e0", X"fa", X"ba", X"41", X"28", X"1b", X"bb", 
    X"ff", X"01", X"1c", X"90", X"00", X"06", X"e0", X"f9", 
    X"a3", X"e0", X"fa", X"eb", X"c3", X"99", X"f9", X"ec", 
    X"9a", X"fa", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e9", X"12", X"17", X"7d", X"a3", X"ea", X"12", X"17", 
    X"7d", X"90", X"05", X"8f", X"e4", X"f0", X"90", X"05", 
    X"8f", X"e0", X"fa", X"70", X"c9", X"22", X"af", X"f0", 
    X"ae", X"83", X"e5", X"82", X"90", X"05", X"90", X"f0", 
    X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"90", X"00", 
    X"00", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"ed", X"4e", X"60", X"33", X"90", X"05", X"90", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"22", 
    X"4f", X"fd", X"a3", X"12", X"22", X"4f", X"fe", X"a3", 
    X"12", X"22", X"4f", X"ff", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"ed", X"12", X"17", X"7d", X"a3", X"ee", 
    X"12", X"17", X"7d", X"a3", X"ef", X"12", X"17", X"7d", 
    X"90", X"00", X"06", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"90", X"00", X"00", X"e0", X"fb", X"a3", X"e0", X"fc", 
    X"a3", X"e0", X"fd", X"74", X"05", X"2b", X"fb", X"e4", 
    X"3c", X"fc", X"90", X"05", X"97", X"ee", X"f0", X"a3", 
    X"ef", X"f0", X"90", X"05", X"99", X"eb", X"f0", X"a3", 
    X"ec", X"f0", X"a3", X"ed", X"f0", X"90", X"00", X"0a", 
    X"02", X"10", X"24", X"90", X"00", X"0a", X"e0", X"ff", 
    X"e4", X"bf", X"41", X"01", X"04", X"ff", X"33", X"95", 
    X"e0", X"fe", X"90", X"00", X"08", X"e0", X"fc", X"a3", 
    X"e0", X"fd", X"90", X"00", X"08", X"ec", X"4f", X"f0", 
    X"ed", X"4e", X"a3", X"f0", X"90", X"00", X"0b", X"74", 
    X"42", X"f0", X"22", X"90", X"00", X"0a", X"74", X"41", 
    X"f0", X"90", X"00", X"08", X"e4", X"f0", X"a3", X"f0", 
    X"22", X"e5", X"82", X"90", X"05", X"96", X"f0", X"90", 
    X"05", X"93", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"90", X"05", X"96", X"e0", X"fc", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"17", X"7d", 
    X"8c", X"82", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"c0", X"04", X"12", X"13", X"74", X"e5", X"82", X"85", 
    X"83", X"f0", X"d0", X"04", X"d0", X"05", X"d0", X"06", 
    X"d0", X"07", X"45", X"f0", X"70", X"0b", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"74", X"03", X"12", X"17", 
    X"7d", X"ec", X"fb", X"24", X"fb", X"40", X"64", X"eb", 
    X"2b", X"2b", X"90", X"0f", X"c6", X"73", X"02", X"0f", 
    X"d5", X"02", X"0f", X"df", X"02", X"10", X"0c", X"02", 
    X"10", X"17", X"02", X"10", X"18", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"e4", X"02", X"17", X"7d", X"90", 
    X"00", X"06", X"e0", X"fb", X"a3", X"e0", X"fc", X"c3", 
    X"74", X"64", X"9b", X"e4", X"64", X"80", X"8c", X"f0", 
    X"63", X"f0", X"80", X"95", X"f0", X"50", X"0a", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"e4", X"02", X"17", 
    X"7d", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", 
    X"03", X"02", X"17", X"7d", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"74", X"01", X"02", X"17", X"7d", X"22", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"02", 
    X"02", X"17", X"7d", X"22", X"af", X"83", X"e5", X"82", 
    X"90", X"05", X"9c", X"f0", X"a3", X"ef", X"f0", X"90", 
    X"05", X"9c", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", 
    X"02", X"2e", X"fe", X"e4", X"3f", X"ff", X"90", X"05", 
    X"99", X"e0", X"fb", X"a3", X"e0", X"fc", X"a3", X"e0", 
    X"fd", X"90", X"05", X"97", X"e0", X"f9", X"a3", X"e0", 
    X"fa", X"ee", X"29", X"fe", X"ef", X"3a", X"ff", X"8b", 
    X"82", X"8c", X"83", X"8d", X"f0", X"ee", X"12", X"17", 
    X"7d", X"a3", X"ef", X"02", X"17", X"7d", X"af", X"f0", 
    X"ae", X"83", X"e5", X"82", X"90", X"05", X"a5", X"f0", 
    X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"90", X"05", 
    X"a1", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"05", 
    X"2e", X"fc", X"e4", X"3f", X"fd", X"90", X"05", X"a5", 
    X"e0", X"f5", X"27", X"a3", X"e0", X"f5", X"28", X"a3", 
    X"e0", X"f5", X"29", X"8c", X"22", X"ed", X"c5", X"22", 
    X"25", X"e0", X"c5", X"22", X"33", X"f5", X"23", X"e5", 
    X"22", X"25", X"27", X"f5", X"24", X"e5", X"23", X"35", 
    X"28", X"f5", X"25", X"85", X"29", X"26", X"90", X"05", 
    X"a3", X"e0", X"f5", X"2a", X"a3", X"e0", X"f5", X"2b", 
    X"85", X"24", X"82", X"85", X"25", X"83", X"85", X"26", 
    X"f0", X"e5", X"2a", X"12", X"17", X"7d", X"a3", X"e5", 
    X"2b", X"12", X"17", X"7d", X"74", X"06", X"2e", X"f9", 
    X"e4", X"3f", X"c9", X"25", X"e0", X"c9", X"33", X"fa", 
    X"e9", X"25", X"27", X"f9", X"ea", X"35", X"28", X"fa", 
    X"ab", X"29", X"89", X"82", X"8a", X"83", X"8b", X"f0", 
    X"e5", X"2a", X"12", X"17", X"7d", X"a3", X"e5", X"2b", 
    X"12", X"17", X"7d", X"74", X"14", X"2e", X"fa", X"e4", 
    X"3f", X"ca", X"25", X"e0", X"ca", X"33", X"fb", X"ea", 
    X"25", X"27", X"fa", X"eb", X"35", X"28", X"f9", X"ab", 
    X"29", X"8a", X"82", X"89", X"83", X"8b", X"f0", X"ec", 
    X"12", X"17", X"7d", X"a3", X"ed", X"12", X"17", X"7d", 
    X"90", X"05", X"9e", X"e0", X"f5", X"30", X"a3", X"e0", 
    X"f5", X"31", X"a3", X"e0", X"f5", X"32", X"90", X"06", 
    X"4c", X"ec", X"f0", X"a3", X"ed", X"f0", X"90", X"00", 
    X"32", X"c0", X"07", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"12", X"17", X"96", X"85", X"82", X"2a", X"85", 
    X"83", X"2b", X"d0", X"04", X"d0", X"05", X"d0", X"06", 
    X"d0", X"07", X"e5", X"2a", X"25", X"30", X"f5", X"27", 
    X"e5", X"2b", X"35", X"31", X"f5", X"28", X"85", X"32", 
    X"29", X"74", X"06", X"2e", X"f5", X"2c", X"e4", X"3f", 
    X"f5", X"2d", X"8c", X"2e", X"8d", X"2f", X"c3", X"e5", 
    X"2c", X"95", X"2e", X"e5", X"2d", X"64", X"80", X"85", 
    X"2f", X"f0", X"63", X"f0", X"80", X"95", X"f0", X"40", 
    X"2c", X"e5", X"2e", X"25", X"2e", X"f8", X"e5", X"2f", 
    X"33", X"fb", X"e8", X"25", X"27", X"f8", X"eb", X"35", 
    X"28", X"fb", X"aa", X"29", X"88", X"82", X"8b", X"83", 
    X"8a", X"f0", X"ec", X"12", X"17", X"7d", X"a3", X"ed", 
    X"12", X"17", X"7d", X"05", X"2e", X"e4", X"b5", X"2e", 
    X"c5", X"05", X"2f", X"80", X"c1", X"e5", X"2a", X"25", 
    X"30", X"f8", X"e5", X"2b", X"35", X"31", X"fa", X"ab", 
    X"32", X"1c", X"ec", X"2c", X"28", X"f8", X"e4", X"3a", 
    X"fa", X"88", X"82", X"8a", X"83", X"8b", X"f0", X"12", 
    X"22", X"4f", X"fc", X"a3", X"12", X"22", X"4f", X"fd", 
    X"0c", X"bc", X"00", X"01", X"0d", X"88", X"82", X"8a", 
    X"83", X"8b", X"f0", X"ec", X"12", X"17", X"7d", X"a3", 
    X"ed", X"12", X"17", X"7d", X"90", X"06", X"4c", X"74", 
    X"0f", X"2e", X"f0", X"e4", X"3f", X"a3", X"f0", X"90", 
    X"00", X"32", X"12", X"17", X"96", X"ae", X"82", X"af", 
    X"83", X"ee", X"25", X"30", X"fe", X"ef", X"35", X"31", 
    X"ff", X"ad", X"32", X"e5", X"22", X"2e", X"fe", X"e5", 
    X"23", X"3f", X"ff", X"85", X"24", X"82", X"85", X"25", 
    X"83", X"85", X"26", X"f0", X"12", X"22", X"4f", X"fb", 
    X"a3", X"12", X"22", X"4f", X"fc", X"8e", X"82", X"8f", 
    X"83", X"8d", X"f0", X"eb", X"12", X"17", X"7d", X"a3", 
    X"ec", X"12", X"17", X"7d", X"90", X"00", X"06", X"74", 
    X"05", X"f0", X"a3", X"e4", X"f0", X"22", X"e5", X"82", 
    X"90", X"05", X"a9", X"f0", X"ff", X"90", X"05", X"a8", 
    X"e0", X"fe", X"ef", X"b5", X"06", X"02", X"80", X"04", 
    X"75", X"82", X"00", X"22", X"90", X"00", X"0a", X"ef", 
    X"f0", X"75", X"82", X"01", X"22", X"af", X"f0", X"ae", 
    X"83", X"e5", X"82", X"90", X"05", X"ad", X"f0", X"a3", 
    X"ee", X"f0", X"a3", X"ef", X"f0", X"90", X"05", X"ad", 
    X"e0", X"f5", X"33", X"a3", X"e0", X"f5", X"34", X"a3", 
    X"e0", X"f5", X"35", X"90", X"05", X"aa", X"e0", X"fa", 
    X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", X"78", X"02", 
    X"79", X"00", X"c3", X"74", X"02", X"98", X"e4", X"64", 
    X"80", X"89", X"f0", X"63", X"f0", X"80", X"95", X"f0", 
    X"40", X"62", X"e8", X"25", X"33", X"fd", X"e9", X"35", 
    X"34", X"fe", X"af", X"35", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"22", X"4f", X"fd", X"74", X"01", 
    X"28", X"fe", X"e4", X"39", X"ff", X"c0", X"00", X"c0", 
    X"01", X"ee", X"2a", X"fe", X"ef", X"3b", X"f9", X"8c", 
    X"07", X"8e", X"82", X"89", X"83", X"8f", X"f0", X"12", 
    X"22", X"4f", X"90", X"05", X"a8", X"f0", X"8d", X"82", 
    X"c0", X"04", X"c0", X"03", X"c0", X"02", X"c0", X"01", 
    X"c0", X"00", X"12", X"12", X"2e", X"e5", X"82", X"d0", 
    X"00", X"d0", X"01", X"d0", X"02", X"d0", X"03", X"d0", 
    X"04", X"d0", X"01", X"d0", X"00", X"70", X"9b", X"90", 
    X"05", X"b2", X"74", X"41", X"f0", X"08", X"b8", X"00", 
    X"91", X"09", X"80", X"8e", X"90", X"05", X"b0", X"e8", 
    X"f0", X"a3", X"e9", X"f0", X"90", X"05", X"b2", X"e0", 
    X"ff", X"c3", X"64", X"80", X"94", X"d7", X"40", X"10", 
    X"ef", X"64", X"80", X"94", X"da", X"50", X"09", X"90", 
    X"05", X"b0", X"74", X"07", X"f0", X"a3", X"e4", X"f0", 
    X"bf", X"52", X"04", X"90", X"00", X"01", X"22", X"90", 
    X"05", X"ad", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"90", X"06", X"4e", X"ea", X"f0", X"a3", 
    X"eb", X"f0", X"a3", X"ec", X"f0", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"17", X"b6", X"ae", X"82", 
    X"af", X"83", X"c3", X"e4", X"9e", X"e4", X"64", X"80", 
    X"8f", X"f0", X"63", X"f0", X"80", X"95", X"f0", X"50", 
    X"27", X"90", X"05", X"b0", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"90", X"05", X"b0", X"74", X"07", X"2e", X"f0", 
    X"e4", X"3f", X"a3", X"f0", X"90", X"05", X"b0", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"90", X"00", X"06", X"ee", 
    X"f0", X"a3", X"ef", X"f0", X"90", X"00", X"01", X"22", 
    X"90", X"00", X"00", X"22", X"e5", X"82", X"90", X"05", 
    X"b3", X"f0", X"ff", X"bf", X"02", X"04", X"90", X"00", 
    X"01", X"22", X"90", X"00", X"00", X"22", X"af", X"83", 
    X"e5", X"82", X"90", X"05", X"b4", X"f0", X"a3", X"ef", 
    X"f0", X"90", X"06", X"1a", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"90", X"06", X"1d", X"ed", 
    X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"90", 
    X"05", X"b4", X"e0", X"fb", X"a3", X"e0", X"fc", X"53", 
    X"03", X"fc", X"90", X"05", X"b4", X"74", X"04", X"2b", 
    X"f0", X"e4", X"3c", X"a3", X"f0", X"90", X"05", X"b4", 
    X"e0", X"fb", X"a3", X"e0", X"fc", X"90", X"06", X"1a", 
    X"eb", X"2d", X"f0", X"ec", X"3e", X"a3", X"f0", X"a3", 
    X"ef", X"f0", X"90", X"06", X"1d", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"22", X"90", X"00", X"00", X"22", 
    X"90", X"00", X"01", X"75", X"f0", X"00", X"22", X"90", 
    X"00", X"00", X"22", X"c0", X"15", X"85", X"81", X"15", 
    X"e5", X"15", X"24", X"fb", X"ff", X"1f", X"1f", X"1f", 
    X"8f", X"01", X"87", X"05", X"09", X"87", X"06", X"09", 
    X"87", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"74", X"30", X"12", X"17", X"7d", X"a3", X"74", X"75", 
    X"12", X"17", X"7d", X"90", X"00", X"00", X"d0", X"15", 
    X"22", X"90", X"06", X"23", X"e4", X"f0", X"a3", X"f0", 
    X"a3", X"f0", X"a3", X"f0", X"90", X"c3", X"50", X"12", 
    X"14", X"c7", X"75", X"82", X"01", X"12", X"15", X"42", 
    X"75", X"82", X"01", X"12", X"14", X"bb", X"75", X"82", 
    X"01", X"02", X"14", X"f1", X"12", X"14", X"fd", X"ae", 
    X"82", X"af", X"83", X"7d", X"00", X"7c", X"00", X"90", 
    X"06", X"37", X"74", X"32", X"f0", X"a3", X"e4", X"f0", 
    X"a3", X"f0", X"a3", X"f0", X"8e", X"82", X"8f", X"83", 
    X"8d", X"f0", X"ec", X"12", X"15", X"fe", X"ac", X"82", 
    X"ad", X"83", X"ae", X"f0", X"ff", X"90", X"06", X"23", 
    X"e0", X"f8", X"a3", X"e0", X"f9", X"a3", X"e0", X"fa", 
    X"a3", X"e0", X"fb", X"90", X"06", X"54", X"e8", X"f0", 
    X"a3", X"e9", X"f0", X"a3", X"ea", X"f0", X"a3", X"eb", 
    X"f0", X"90", X"03", X"e8", X"e4", X"f5", X"f0", X"c0", 
    X"07", X"c0", X"06", X"c0", X"05", X"c0", X"04", X"12", 
    X"18", X"4a", X"a8", X"82", X"a9", X"83", X"aa", X"f0", 
    X"fb", X"d0", X"04", X"d0", X"05", X"d0", X"06", X"d0", 
    X"07", X"e8", X"2c", X"fc", X"e9", X"3d", X"fd", X"ea", 
    X"3e", X"fe", X"eb", X"3f", X"8c", X"82", X"8d", X"83", 
    X"8e", X"f0", X"22", X"e5", X"82", X"90", X"06", X"27", 
    X"f0", X"13", X"92", X"00", X"92", X"af", X"22", X"af", 
    X"83", X"e5", X"82", X"90", X"06", X"28", X"f0", X"a3", 
    X"ef", X"f0", X"90", X"06", X"28", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"be", X"ff", X"05", X"bf", X"ff", X"02", 
    X"80", X"0a", X"8f", X"8f", X"7f", X"00", X"8e", X"8e", 
    X"d2", X"8c", X"80", X"02", X"c2", X"8c", X"d2", X"88", 
    X"22", X"e5", X"82", X"90", X"06", X"2a", X"f0", X"13", 
    X"92", X"01", X"92", X"8d", X"22", X"90", X"06", X"2b", 
    X"e5", X"8d", X"f0", X"90", X"06", X"2c", X"e5", X"8c", 
    X"f0", X"90", X"06", X"2d", X"e5", X"8c", X"f0", X"90", 
    X"06", X"2c", X"e0", X"ff", X"90", X"06", X"2d", X"e0", 
    X"fe", X"ef", X"b5", X"06", X"02", X"80", X"0c", X"90", 
    X"06", X"2b", X"e5", X"8d", X"f0", X"90", X"06", X"2c", 
    X"e5", X"8c", X"f0", X"90", X"06", X"2b", X"e0", X"fe", 
    X"7f", X"00", X"90", X"06", X"2c", X"e0", X"7c", X"00", 
    X"42", X"07", X"ec", X"42", X"06", X"8f", X"82", X"8e", 
    X"83", X"22", X"e5", X"82", X"90", X"06", X"2e", X"f0", 
    X"13", X"92", X"02", X"92", X"a9", X"22", X"c0", X"e0", 
    X"c0", X"82", X"c0", X"83", X"c0", X"07", X"c0", X"d0", 
    X"75", X"d0", X"00", X"d2", X"88", X"90", X"06", X"2f", 
    X"e0", X"ff", X"8f", X"90", X"90", X"06", X"2f", X"ef", 
    X"04", X"f0", X"90", X"06", X"23", X"e0", X"24", X"01", 
    X"f0", X"a3", X"e0", X"34", X"00", X"f0", X"a3", X"e0", 
    X"34", X"00", X"f0", X"a3", X"e0", X"34", X"00", X"f0", 
    X"d0", X"d0", X"d0", X"07", X"d0", X"83", X"d0", X"82", 
    X"d0", X"e0", X"32", X"e5", X"82", X"90", X"06", X"30", 
    X"f0", X"30", X"9c", X"fd", X"90", X"06", X"30", X"e0", 
    X"ff", X"8f", X"99", X"bf", X"0a", X"06", X"30", X"9c", 
    X"fd", X"75", X"99", X"0d", X"22", X"af", X"f0", X"ae", 
    X"83", X"e5", X"82", X"90", X"06", X"34", X"f0", X"a3", 
    X"ee", X"f0", X"a3", X"ef", X"f0", X"90", X"06", X"34", 
    X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"90", X"06", X"31", X"e0", X"fa", X"a3", X"e0", X"fb", 
    X"a3", X"e0", X"fc", X"8d", X"36", X"8e", X"37", X"8f", 
    X"38", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", 
    X"22", X"4f", X"f9", X"a3", X"aa", X"82", X"ab", X"83", 
    X"85", X"36", X"82", X"85", X"37", X"83", X"85", X"38", 
    X"f0", X"e9", X"12", X"17", X"7d", X"a3", X"85", X"82", 
    X"36", X"85", X"83", X"37", X"e9", X"70", X"da", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"22", X"af", X"82", 
    X"ae", X"83", X"ad", X"f0", X"fc", X"90", X"06", X"3b", 
    X"ef", X"f0", X"a3", X"ee", X"f0", X"a3", X"ed", X"f0", 
    X"a3", X"ec", X"f0", X"90", X"06", X"3f", X"e4", X"f0", 
    X"a3", X"f0", X"a3", X"f0", X"a3", X"f0", X"90", X"06", 
    X"37", X"e0", X"fc", X"a3", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"75", X"36", X"20", X"90", 
    X"06", X"3b", X"e0", X"f8", X"a3", X"e0", X"f9", X"a3", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"33", X"92", X"03", 
    X"e8", X"28", X"f8", X"e9", X"33", X"f9", X"ea", X"33", 
    X"fa", X"eb", X"33", X"fb", X"90", X"06", X"3b", X"e8", 
    X"f0", X"a3", X"e9", X"f0", X"a3", X"ea", X"f0", X"a3", 
    X"eb", X"f0", X"90", X"06", X"3f", X"e0", X"f8", X"a3", 
    X"e0", X"f9", X"a3", X"e0", X"fa", X"a3", X"e0", X"fb", 
    X"e8", X"28", X"f8", X"e9", X"33", X"f9", X"ea", X"33", 
    X"fa", X"eb", X"33", X"fb", X"90", X"06", X"3f", X"e8", 
    X"f0", X"a3", X"e9", X"f0", X"a3", X"ea", X"f0", X"a3", 
    X"eb", X"f0", X"30", X"03", X"1e", X"90", X"06", X"3f", 
    X"e0", X"f8", X"a3", X"e0", X"f9", X"a3", X"e0", X"fa", 
    X"a3", X"e0", X"fb", X"90", X"06", X"3f", X"74", X"01", 
    X"48", X"f0", X"a3", X"e9", X"f0", X"a3", X"ea", X"f0", 
    X"a3", X"eb", X"f0", X"90", X"06", X"3f", X"e0", X"f8", 
    X"a3", X"e0", X"f9", X"a3", X"e0", X"fa", X"a3", X"e0", 
    X"fb", X"c3", X"e8", X"9c", X"e9", X"9d", X"ea", X"9e", 
    X"eb", X"9f", X"40", X"31", X"90", X"06", X"3f", X"e8", 
    X"c3", X"9c", X"f0", X"e9", X"9d", X"a3", X"f0", X"ea", 
    X"9e", X"a3", X"f0", X"eb", X"9f", X"a3", X"f0", X"90", 
    X"06", X"3b", X"e0", X"f8", X"a3", X"e0", X"f9", X"a3", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"90", X"06", X"3b", 
    X"74", X"01", X"48", X"f0", X"a3", X"e9", X"f0", X"a3", 
    X"ea", X"f0", X"a3", X"eb", X"f0", X"d5", X"36", X"02", 
    X"80", X"03", X"02", X"16", X"2f", X"90", X"06", X"3b", 
    X"e0", X"fc", X"a3", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"8c", X"82", X"8d", X"83", X"8e", X"f0", 
    X"22", X"af", X"f0", X"ae", X"83", X"e5", X"82", X"90", 
    X"06", X"48", X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", 
    X"f0", X"90", X"06", X"48", X"e0", X"f5", X"36", X"a3", 
    X"e0", X"f5", X"37", X"a3", X"e0", X"f5", X"38", X"aa", 
    X"36", X"ab", X"37", X"ac", X"38", X"90", X"06", X"43", 
    X"e0", X"f8", X"a3", X"e0", X"f9", X"a3", X"e0", X"ff", 
    X"90", X"06", X"46", X"e0", X"f5", X"39", X"a3", X"e0", 
    X"f5", X"3a", X"ad", X"39", X"ae", X"3a", X"15", X"39", 
    X"74", X"ff", X"b5", X"39", X"02", X"15", X"3a", X"ed", 
    X"4e", X"60", X"20", X"88", X"82", X"89", X"83", X"8f", 
    X"f0", X"12", X"22", X"4f", X"fe", X"a3", X"a8", X"82", 
    X"a9", X"83", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"ee", X"12", X"17", X"7d", X"a3", X"aa", X"82", X"ab", 
    X"83", X"80", X"cf", X"85", X"36", X"82", X"85", X"37", 
    X"83", X"85", X"38", X"f0", X"22", X"20", X"f7", X"10", 
    X"30", X"f6", X"11", X"88", X"83", X"a8", X"82", X"20", 
    X"f5", X"07", X"f6", X"a8", X"83", X"75", X"83", X"00", 
    X"22", X"f2", X"80", X"f7", X"f0", X"22", X"aa", X"83", 
    X"ab", X"82", X"8b", X"f0", X"90", X"06", X"4c", X"e0", 
    X"a4", X"f8", X"a9", X"f0", X"8a", X"f0", X"e0", X"a4", 
    X"29", X"f9", X"8b", X"f0", X"a3", X"e0", X"a4", X"29", 
    X"f5", X"83", X"88", X"82", X"22", X"22", X"af", X"f0", 
    X"ae", X"83", X"e5", X"82", X"90", X"06", X"51", X"f0", 
    X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"90", X"06", 
    X"51", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"90", X"06", X"4e", X"e0", X"f5", X"36", X"a3", 
    X"e0", X"f5", X"37", X"a3", X"e0", X"f5", X"38", X"8d", 
    X"00", X"8e", X"01", X"8f", X"04", X"88", X"82", X"89", 
    X"83", X"8c", X"f0", X"12", X"22", X"4f", X"f8", X"7c", 
    X"00", X"a9", X"36", X"aa", X"37", X"ab", X"38", X"89", 
    X"82", X"8a", X"83", X"8b", X"f0", X"12", X"22", X"4f", 
    X"f9", X"7b", X"00", X"e8", X"c3", X"99", X"f8", X"ec", 
    X"9b", X"fc", X"88", X"02", X"8c", X"03", X"e8", X"4c", 
    X"70", X"28", X"85", X"36", X"82", X"85", X"37", X"83", 
    X"85", X"38", X"f0", X"12", X"22", X"4f", X"60", X"1a", 
    X"0d", X"bd", X"00", X"01", X"0e", X"90", X"06", X"51", 
    X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", 
    X"05", X"36", X"e4", X"b5", X"36", X"a9", X"05", X"37", 
    X"80", X"a5", X"90", X"06", X"51", X"ed", X"f0", X"a3", 
    X"ee", X"f0", X"a3", X"ef", X"f0", X"8a", X"82", X"8b", 
    X"83", X"22", X"a8", X"82", X"a9", X"83", X"aa", X"f0", 
    X"fb", X"88", X"f0", X"90", X"06", X"54", X"e0", X"a4", 
    X"fc", X"ad", X"f0", X"89", X"f0", X"e0", X"a4", X"2d", 
    X"fd", X"e4", X"35", X"f0", X"fe", X"88", X"f0", X"a3", 
    X"e0", X"a4", X"2d", X"fd", X"e5", X"f0", X"3e", X"fe", 
    X"e4", X"33", X"ff", X"89", X"f0", X"e0", X"a4", X"2e", 
    X"fe", X"e5", X"f0", X"3f", X"ff", X"88", X"f0", X"a3", 
    X"e0", X"a4", X"2e", X"fe", X"e5", X"f0", X"3f", X"ff", 
    X"8a", X"f0", X"90", X"06", X"54", X"e0", X"a4", X"2e", 
    X"fe", X"e5", X"f0", X"3f", X"ff", X"8b", X"f0", X"e0", 
    X"a4", X"2f", X"ff", X"8a", X"f0", X"a3", X"e0", X"a4", 
    X"2f", X"ff", X"89", X"f0", X"a3", X"e0", X"a4", X"2f", 
    X"ff", X"88", X"f0", X"a3", X"e0", X"a4", X"2f", X"8e", 
    X"f0", X"8d", X"83", X"8c", X"82", X"22", X"af", X"83", 
    X"e5", X"82", X"90", X"06", X"5a", X"f0", X"a3", X"ef", 
    X"f0", X"90", X"06", X"5a", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"33", X"e4", X"33", X"fd", X"60", X"09", X"c3", 
    X"e4", X"9e", X"fb", X"e4", X"9f", X"fc", X"80", X"04", 
    X"8e", X"03", X"8f", X"04", X"90", X"06", X"58", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"33", X"e4", X"33", X"fa", 
    X"60", X"09", X"c3", X"e4", X"9e", X"f8", X"e4", X"9f", 
    X"f9", X"80", X"04", X"8e", X"00", X"8f", X"01", X"90", 
    X"06", X"5c", X"e8", X"f0", X"a3", X"e9", X"f0", X"8b", 
    X"82", X"8c", X"83", X"c0", X"05", X"c0", X"02", X"12", 
    X"19", X"27", X"ae", X"82", X"af", X"83", X"d0", X"02", 
    X"d0", X"05", X"ea", X"6d", X"60", X"0c", X"c3", X"e4", 
    X"9e", X"fc", X"e4", X"9f", X"fd", X"8c", X"82", X"8d", 
    X"83", X"22", X"8e", X"82", X"8f", X"83", X"22", X"af", 
    X"83", X"e5", X"82", X"90", X"06", X"5e", X"f0", X"a3", 
    X"ef", X"f0", X"90", X"06", X"60", X"e4", X"f0", X"a3", 
    X"f0", X"90", X"06", X"5c", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"7d", X"10", X"90", X"06", X"5e", X"e0", X"fb", 
    X"a3", X"e0", X"fc", X"33", X"92", X"04", X"ec", X"cb", 
    X"25", X"e0", X"cb", X"33", X"fc", X"90", X"06", X"5e", 
    X"eb", X"f0", X"a3", X"ec", X"f0", X"90", X"06", X"60", 
    X"e0", X"fb", X"a3", X"e0", X"cb", X"25", X"e0", X"cb", 
    X"33", X"fc", X"90", X"06", X"60", X"eb", X"f0", X"a3", 
    X"ec", X"f0", X"30", X"04", X"12", X"90", X"06", X"60", 
    X"e0", X"fb", X"a3", X"e0", X"fc", X"90", X"06", X"60", 
    X"74", X"01", X"4b", X"f0", X"a3", X"ec", X"f0", X"90", 
    X"06", X"60", X"e0", X"fb", X"a3", X"e0", X"fc", X"c3", 
    X"eb", X"9e", X"ec", X"9f", X"40", X"1d", X"90", X"06", 
    X"60", X"eb", X"c3", X"9e", X"f0", X"ec", X"9f", X"a3", 
    X"f0", X"90", X"06", X"5e", X"e0", X"fb", X"a3", X"e0", 
    X"fc", X"90", X"06", X"5e", X"74", X"01", X"4b", X"f0", 
    X"a3", X"ec", X"f0", X"dd", X"8e", X"90", X"06", X"5e", 
    X"e0", X"fe", X"a3", X"e0", X"8e", X"82", X"f5", X"83", 
    X"22", X"c0", X"15", X"85", X"81", X"15", X"12", X"15", 
    X"8b", X"d0", X"15", X"22", X"af", X"f0", X"ae", X"83", 
    X"e5", X"82", X"90", X"06", X"63", X"f0", X"a3", X"ee", 
    X"f0", X"a3", X"ef", X"f0", X"90", X"06", X"63", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"90", 
    X"06", X"62", X"e0", X"fc", X"90", X"06", X"76", X"e4", 
    X"f0", X"a3", X"f0", X"a3", X"f0", X"90", X"06", X"79", 
    X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", 
    X"90", X"06", X"7c", X"ec", X"f0", X"90", X"19", X"c1", 
    X"02", X"1b", X"0e", X"c0", X"15", X"85", X"81", X"15", 
    X"e5", X"15", X"24", X"fb", X"ff", X"90", X"06", X"76", 
    X"e4", X"f0", X"a3", X"f0", X"a3", X"f0", X"e5", X"15", 
    X"24", X"fb", X"f8", X"90", X"06", X"79", X"e6", X"f0", 
    X"08", X"a3", X"e6", X"f0", X"08", X"a3", X"e6", X"f0", 
    X"90", X"06", X"7c", X"ef", X"f0", X"90", X"19", X"c1", 
    X"12", X"1b", X"0e", X"d0", X"15", X"22", X"e5", X"82", 
    X"90", X"06", X"72", X"f0", X"ff", X"90", X"06", X"68", 
    X"e0", X"c0", X"e0", X"a3", X"e0", X"c0", X"e0", X"a3", 
    X"e0", X"c0", X"e0", X"74", X"68", X"c0", X"e0", X"74", 
    X"1a", X"c0", X"e0", X"90", X"06", X"66", X"e0", X"c0", 
    X"e0", X"a3", X"e0", X"c0", X"e0", X"8f", X"82", X"22", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"90", X"06", 
    X"70", X"e0", X"24", X"01", X"f0", X"a3", X"e0", X"34", 
    X"00", X"f0", X"22", X"e5", X"82", X"90", X"06", X"73", 
    X"f0", X"24", X"30", X"ff", X"24", X"c6", X"50", X"0a", 
    X"74", X"07", X"2f", X"ff", X"30", X"05", X"03", X"43", 
    X"07", X"20", X"8f", X"82", X"02", X"1a", X"3e", X"e5", 
    X"82", X"90", X"06", X"74", X"f0", X"ff", X"c4", X"54", 
    X"0f", X"f5", X"82", X"c0", X"07", X"12", X"1a", X"7b", 
    X"d0", X"07", X"53", X"07", X"0f", X"8f", X"82", X"02", 
    X"1a", X"7b", X"e5", X"82", X"90", X"06", X"75", X"f0", 
    X"90", X"06", X"6b", X"e0", X"fc", X"a3", X"e0", X"fd", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"90", X"06", 
    X"6f", X"e0", X"fb", X"90", X"06", X"75", X"e0", X"fa", 
    X"75", X"36", X"20", X"eb", X"2b", X"fb", X"ef", X"23", 
    X"54", X"01", X"f8", X"8b", X"01", X"49", X"fb", X"ec", 
    X"2c", X"fc", X"ed", X"33", X"fd", X"ee", X"33", X"fe", 
    X"ef", X"33", X"ff", X"c3", X"eb", X"9a", X"40", X"07", 
    X"eb", X"c3", X"9a", X"fb", X"43", X"04", X"01", X"d5", 
    X"36", X"d9", X"90", X"06", X"6b", X"ec", X"f0", X"a3", 
    X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", 
    X"90", X"06", X"6f", X"eb", X"f0", X"22", X"af", X"83", 
    X"e5", X"82", X"90", X"06", X"7d", X"f0", X"a3", X"ef", 
    X"f0", X"90", X"06", X"7d", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"90", X"06", X"66", X"ee", X"f0", X"a3", X"ef", 
    X"f0", X"90", X"06", X"76", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"90", X"06", X"68", X"ed", 
    X"f0", X"a3", X"ee", X"f0", X"a3", X"ef", X"f0", X"90", 
    X"06", X"70", X"e4", X"f0", X"a3", X"f0", X"90", X"06", 
    X"79", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"22", X"4f", X"fc", X"90", X"06", X"79", X"74", X"01", 
    X"2d", X"f0", X"e4", X"3e", X"a3", X"f0", X"a3", X"ef", 
    X"f0", X"ec", X"70", X"03", X"02", X"22", X"2b", X"bc", 
    X"25", X"02", X"80", X"03", X"02", X"22", X"23", X"c2", 
    X"06", X"c2", X"07", X"c2", X"08", X"c2", X"09", X"c2", 
    X"0a", X"c2", X"0b", X"c2", X"0c", X"c2", X"0d", X"90", 
    X"06", X"7f", X"e4", X"f0", X"90", X"06", X"80", X"f0", 
    X"90", X"06", X"81", X"74", X"ff", X"f0", X"90", X"06", 
    X"79", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"22", X"4f", X"fb", X"a3", X"ad", X"82", X"ae", X"83", 
    X"90", X"06", X"79", X"ed", X"f0", X"a3", X"ee", X"f0", 
    X"a3", X"ef", X"f0", X"90", X"06", X"83", X"eb", X"f0", 
    X"bb", X"25", X"08", X"8b", X"82", X"12", X"1a", X"3e", 
    X"02", X"1b", X"46", X"8b", X"02", X"ba", X"30", X"00", 
    X"40", X"3c", X"ea", X"24", X"c6", X"40", X"37", X"90", 
    X"06", X"81", X"e0", X"fa", X"ba", X"ff", X"21", X"c0", 
    X"05", X"c0", X"06", X"c0", X"07", X"90", X"06", X"80", 
    X"e0", X"75", X"f0", X"0a", X"a4", X"2b", X"24", X"d0", 
    X"90", X"06", X"80", X"f0", X"d0", X"07", X"d0", X"06", 
    X"d0", X"05", X"70", X"a5", X"d2", X"07", X"80", X"a1", 
    X"ea", X"75", X"f0", X"0a", X"a4", X"2b", X"24", X"d0", 
    X"90", X"06", X"81", X"f0", X"80", X"93", X"90", X"06", 
    X"83", X"e0", X"fb", X"bb", X"2e", X"15", X"90", X"06", 
    X"81", X"e0", X"fa", X"ba", X"ff", X"02", X"80", X"03", 
    X"02", X"1b", X"a1", X"90", X"06", X"81", X"e4", X"f0", 
    X"02", X"1b", X"a1", X"8b", X"02", X"ba", X"61", X"00", 
    X"40", X"10", X"ea", X"24", X"85", X"40", X"0b", X"90", 
    X"06", X"83", X"74", X"df", X"5b", X"f0", X"d2", X"05", 
    X"80", X"02", X"c2", X"05", X"90", X"06", X"83", X"e0", 
    X"fb", X"bb", X"20", X"02", X"80", X"6d", X"bb", X"2b", 
    X"02", X"80", X"63", X"bb", X"2d", X"02", X"80", X"59", 
    X"bb", X"42", X"02", X"80", X"63", X"bb", X"43", X"02", 
    X"80", X"68", X"bb", X"44", X"03", X"02", X"1e", X"aa", 
    X"bb", X"46", X"03", X"02", X"1e", X"cc", X"bb", X"48", 
    X"03", X"02", X"1b", X"a1", X"bb", X"49", X"03", X"02", 
    X"1e", X"aa", X"bb", X"4a", X"03", X"02", X"1b", X"a1", 
    X"bb", X"4c", X"02", X"80", X"40", X"bb", X"4f", X"03", 
    X"02", X"1e", X"b4", X"bb", X"50", X"03", X"02", X"1e", 
    X"16", X"bb", X"53", X"02", X"80", X"70", X"bb", X"54", 
    X"03", X"02", X"1b", X"a1", X"bb", X"55", X"03", X"02", 
    X"1e", X"bc", X"bb", X"58", X"03", X"02", X"1e", X"c4", 
    X"bb", X"5a", X"03", X"02", X"1b", X"a1", X"02", X"1e", 
    X"d0", X"d2", X"06", X"02", X"1b", X"a1", X"d2", X"08", 
    X"02", X"1b", X"a1", X"d2", X"09", X"02", X"1b", X"a1", 
    X"d2", X"0b", X"02", X"1b", X"a1", X"d2", X"0c", X"02", 
    X"1b", X"a1", X"30", X"0b", X"14", X"90", X"06", X"7c", 
    X"e0", X"ff", X"1f", X"90", X"06", X"7c", X"ef", X"f0", 
    X"8f", X"01", X"90", X"06", X"83", X"e7", X"f0", X"80", 
    X"19", X"90", X"06", X"7c", X"e0", X"ff", X"1f", X"1f", 
    X"90", X"06", X"7c", X"ef", X"f0", X"8f", X"01", X"87", 
    X"06", X"09", X"87", X"07", X"19", X"90", X"06", X"83", 
    X"ee", X"f0", X"90", X"06", X"83", X"e0", X"f5", X"82", 
    X"12", X"1a", X"3e", X"02", X"1e", X"dc", X"90", X"06", 
    X"7c", X"e0", X"ff", X"1f", X"1f", X"1f", X"90", X"06", 
    X"7c", X"ef", X"f0", X"8f", X"01", X"87", X"05", X"09", 
    X"87", X"06", X"09", X"87", X"07", X"19", X"19", X"90", 
    X"06", X"6b", X"ed", X"f0", X"a3", X"ee", X"f0", X"a3", 
    X"ef", X"f0", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"22", X"37", X"ae", X"82", X"90", X"06", X"81", 
    X"e0", X"ff", X"bf", X"ff", X"05", X"90", X"06", X"81", 
    X"ee", X"f0", X"20", X"06", X"36", X"90", X"06", X"80", 
    X"e0", X"ff", X"c3", X"ee", X"9f", X"50", X"2c", X"90", 
    X"06", X"80", X"ef", X"c3", X"9e", X"f0", X"90", X"06", 
    X"80", X"e0", X"ff", X"8f", X"05", X"1f", X"90", X"06", 
    X"80", X"ef", X"f0", X"ed", X"60", X"10", X"75", X"82", 
    X"20", X"c0", X"07", X"c0", X"06", X"12", X"1a", X"3e", 
    X"d0", X"06", X"d0", X"07", X"80", X"e5", X"90", X"06", 
    X"80", X"ef", X"f0", X"90", X"06", X"81", X"e0", X"ff", 
    X"c0", X"06", X"90", X"06", X"6b", X"e0", X"fa", X"a3", 
    X"e0", X"fd", X"a3", X"e0", X"fe", X"8a", X"82", X"8d", 
    X"83", X"8e", X"f0", X"12", X"22", X"4f", X"f5", X"16", 
    X"d0", X"06", X"e5", X"16", X"60", X"3f", X"8f", X"05", 
    X"1f", X"c3", X"e4", X"64", X"80", X"8d", X"f0", X"63", 
    X"f0", X"80", X"95", X"f0", X"50", X"2f", X"c0", X"06", 
    X"85", X"16", X"82", X"c0", X"07", X"c0", X"06", X"12", 
    X"1a", X"3e", X"d0", X"06", X"d0", X"07", X"90", X"06", 
    X"6b", X"e0", X"fa", X"a3", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"0a", X"ba", X"00", X"01", X"0d", X"90", X"06", 
    X"6b", X"ea", X"f0", X"a3", X"ed", X"f0", X"a3", X"ee", 
    X"f0", X"d0", X"06", X"80", X"a3", X"20", X"06", X"03", 
    X"02", X"1e", X"dc", X"90", X"06", X"80", X"e0", X"ff", 
    X"c3", X"ee", X"9f", X"40", X"03", X"02", X"1e", X"dc", 
    X"90", X"06", X"80", X"ef", X"c3", X"9e", X"f0", X"90", 
    X"06", X"80", X"e0", X"ff", X"8f", X"06", X"1f", X"90", 
    X"06", X"80", X"ef", X"f0", X"ee", X"70", X"03", X"02", 
    X"1e", X"d7", X"75", X"82", X"20", X"c0", X"07", X"12", 
    X"1a", X"3e", X"d0", X"07", X"80", X"e6", X"90", X"06", 
    X"7c", X"e0", X"fe", X"1e", X"1e", X"1e", X"90", X"06", 
    X"7c", X"ee", X"f0", X"8e", X"01", X"87", X"02", X"09", 
    X"87", X"05", X"09", X"87", X"06", X"19", X"19", X"90", 
    X"06", X"6b", X"ea", X"f0", X"a3", X"ed", X"f0", X"a3", 
    X"ee", X"f0", X"90", X"06", X"6d", X"e0", X"fe", X"be", 
    X"80", X"00", X"40", X"08", X"90", X"06", X"83", X"74", 
    X"43", X"f0", X"80", X"20", X"be", X"60", X"00", X"40", 
    X"08", X"90", X"06", X"83", X"74", X"50", X"f0", X"80", 
    X"13", X"be", X"40", X"00", X"40", X"08", X"90", X"06", 
    X"83", X"74", X"49", X"f0", X"80", X"06", X"90", X"06", 
    X"83", X"74", X"58", X"f0", X"90", X"06", X"83", X"e0", 
    X"fe", X"f5", X"82", X"c0", X"06", X"12", X"1a", X"3e", 
    X"75", X"82", X"3a", X"12", X"1a", X"3e", X"75", X"82", 
    X"30", X"12", X"1a", X"3e", X"75", X"82", X"78", X"12", 
    X"1a", X"3e", X"d0", X"06", X"be", X"49", X"02", X"80", 
    X"0e", X"be", X"50", X"02", X"80", X"09", X"90", X"06", 
    X"6c", X"e0", X"f5", X"82", X"12", X"1a", X"97", X"90", 
    X"06", X"6b", X"e0", X"f5", X"82", X"12", X"1a", X"97", 
    X"80", X"32", X"d2", X"0a", X"90", X"06", X"7f", X"74", 
    X"0a", X"f0", X"80", X"28", X"90", X"06", X"7f", X"74", 
    X"08", X"f0", X"80", X"20", X"90", X"06", X"7f", X"74", 
    X"0a", X"f0", X"80", X"18", X"90", X"06", X"7f", X"74", 
    X"10", X"f0", X"80", X"10", X"d2", X"0d", X"80", X"0c", 
    X"8b", X"82", X"12", X"1a", X"3e", X"80", X"05", X"90", 
    X"06", X"80", X"ef", X"f0", X"30", X"0d", X"77", X"90", 
    X"06", X"7c", X"e0", X"ff", X"1f", X"1f", X"1f", X"1f", 
    X"90", X"06", X"7c", X"ef", X"f0", X"8f", X"01", X"87", 
    X"03", X"09", X"87", X"05", X"09", X"87", X"06", X"09", 
    X"87", X"07", X"19", X"19", X"19", X"90", X"06", X"6b", 
    X"eb", X"f0", X"a3", X"ed", X"f0", X"a3", X"ee", X"f0", 
    X"a3", X"ef", X"f0", X"90", X"06", X"6b", X"74", X"57", 
    X"f0", X"a3", X"74", X"27", X"f0", X"a3", X"74", X"80", 
    X"f0", X"90", X"06", X"6b", X"e0", X"f5", X"17", X"a3", 
    X"e0", X"f5", X"18", X"a3", X"e0", X"f5", X"19", X"74", 
    X"01", X"25", X"17", X"fa", X"e4", X"35", X"18", X"fb", 
    X"af", X"19", X"90", X"06", X"6b", X"ea", X"f0", X"a3", 
    X"eb", X"f0", X"a3", X"ef", X"f0", X"85", X"17", X"82", 
    X"85", X"18", X"83", X"85", X"19", X"f0", X"12", X"22", 
    X"4f", X"ff", X"70", X"03", X"02", X"1b", X"46", X"8f", 
    X"82", X"12", X"1a", X"3e", X"80", X"c3", X"90", X"06", 
    X"7f", X"e0", X"f5", X"17", X"70", X"03", X"02", X"1b", 
    X"46", X"90", X"06", X"8a", X"74", X"89", X"f0", X"a3", 
    X"74", X"06", X"f0", X"30", X"0b", X"4a", X"90", X"06", 
    X"7c", X"e0", X"fe", X"1e", X"90", X"06", X"7c", X"ee", 
    X"f0", X"8e", X"01", X"e7", X"fe", X"33", X"95", X"e0", 
    X"fd", X"fb", X"fa", X"90", X"06", X"6b", X"ee", X"f0", 
    X"a3", X"ed", X"f0", X"a3", X"eb", X"f0", X"a3", X"ea", 
    X"f0", X"30", X"0a", X"03", X"02", X"20", X"32", X"90", 
    X"06", X"6b", X"e0", X"fa", X"a3", X"e0", X"a3", X"e0", 
    X"a3", X"e0", X"7b", X"00", X"7d", X"00", X"7e", X"00", 
    X"90", X"06", X"6b", X"ea", X"f0", X"a3", X"eb", X"f0", 
    X"a3", X"ed", X"f0", X"a3", X"ee", X"f0", X"80", X"7a", 
    X"30", X"0c", X"2e", X"90", X"06", X"7c", X"e0", X"fe", 
    X"1e", X"1e", X"1e", X"1e", X"90", X"06", X"7c", X"ee", 
    X"f0", X"8e", X"01", X"87", X"02", X"09", X"87", X"03", 
    X"09", X"87", X"05", X"09", X"87", X"06", X"19", X"19", 
    X"19", X"90", X"06", X"6b", X"ea", X"f0", X"a3", X"eb", 
    X"f0", X"a3", X"ed", X"f0", X"a3", X"ee", X"f0", X"80", 
    X"49", X"90", X"06", X"7c", X"e0", X"fe", X"1e", X"1e", 
    X"90", X"06", X"7c", X"ee", X"f0", X"8e", X"01", X"87", 
    X"05", X"09", X"87", X"06", X"19", X"ee", X"33", X"95", 
    X"e0", X"fb", X"fa", X"90", X"06", X"6b", X"ed", X"f0", 
    X"a3", X"ee", X"f0", X"a3", X"eb", X"f0", X"a3", X"ea", 
    X"f0", X"20", X"0a", X"1e", X"90", X"06", X"6b", X"e0", 
    X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"a3", X"e0", 
    X"7d", X"00", X"7e", X"00", X"90", X"06", X"6b", X"ea", 
    X"f0", X"a3", X"eb", X"f0", X"a3", X"ed", X"f0", X"a3", 
    X"ee", X"f0", X"30", X"0a", X"30", X"90", X"06", X"6b", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"fd", 
    X"a3", X"e0", X"fe", X"30", X"e7", X"1d", X"c3", X"e4", 
    X"9a", X"fa", X"e4", X"9b", X"fb", X"e4", X"9d", X"fd", 
    X"e4", X"9e", X"fe", X"90", X"06", X"6b", X"ea", X"f0", 
    X"a3", X"eb", X"f0", X"a3", X"ed", X"f0", X"a3", X"ee", 
    X"f0", X"80", X"02", X"c2", X"0a", X"d2", X"0e", X"75", 
    X"1a", X"89", X"75", X"1b", X"06", X"75", X"16", X"00", 
    X"90", X"06", X"6f", X"e4", X"f0", X"85", X"17", X"82", 
    X"12", X"1a", X"b2", X"20", X"0e", X"2d", X"90", X"06", 
    X"6f", X"e0", X"c4", X"fa", X"85", X"1a", X"82", X"85", 
    X"1b", X"83", X"e0", X"ff", X"42", X"02", X"85", X"1a", 
    X"82", X"85", X"1b", X"83", X"ea", X"f0", X"15", X"1a", 
    X"74", X"ff", X"b5", X"1a", X"02", X"15", X"1b", X"90", 
    X"06", X"8a", X"e5", X"1a", X"f0", X"a3", X"e5", X"1b", 
    X"f0", X"80", X"0c", X"90", X"06", X"6f", X"e0", X"fa", 
    X"85", X"1a", X"82", X"85", X"1b", X"83", X"f0", X"05", 
    X"16", X"90", X"06", X"82", X"e5", X"16", X"f0", X"b2", 
    X"0e", X"90", X"06", X"6b", X"e0", X"fa", X"a3", X"e0", 
    X"fb", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"ea", 
    X"4b", X"4e", X"4f", X"70", X"9b", X"90", X"06", X"8a", 
    X"e5", X"1a", X"f0", X"a3", X"e5", X"1b", X"f0", X"90", 
    X"06", X"82", X"e5", X"16", X"f0", X"90", X"06", X"80", 
    X"e0", X"ff", X"70", X"06", X"90", X"06", X"80", X"74", 
    X"01", X"f0", X"20", X"07", X"27", X"20", X"06", X"24", 
    X"e5", X"16", X"04", X"ff", X"90", X"06", X"80", X"e0", 
    X"fe", X"c3", X"ef", X"9e", X"50", X"11", X"75", X"82", 
    X"20", X"c0", X"07", X"c0", X"06", X"12", X"1a", X"3e", 
    X"d0", X"06", X"d0", X"07", X"1e", X"80", X"ea", X"90", 
    X"06", X"80", X"ee", X"f0", X"30", X"0a", X"11", X"75", 
    X"82", X"2d", X"12", X"1a", X"3e", X"90", X"06", X"80", 
    X"e0", X"14", X"90", X"06", X"80", X"f0", X"80", X"2d", 
    X"90", X"06", X"82", X"e0", X"ff", X"60", X"26", X"30", 
    X"08", X"11", X"75", X"82", X"2b", X"12", X"1a", X"3e", 
    X"90", X"06", X"80", X"e0", X"14", X"90", X"06", X"80", 
    X"f0", X"80", X"12", X"30", X"09", X"0f", X"75", X"82", 
    X"20", X"12", X"1a", X"3e", X"90", X"06", X"80", X"e0", 
    X"14", X"90", X"06", X"80", X"f0", X"20", X"06", X"2f", 
    X"90", X"06", X"82", X"e0", X"ff", X"90", X"06", X"80", 
    X"e0", X"fe", X"8e", X"05", X"1e", X"90", X"06", X"80", 
    X"ee", X"f0", X"c3", X"ef", X"9d", X"50", X"36", X"30", 
    X"07", X"04", X"7d", X"30", X"80", X"02", X"7d", X"20", 
    X"8d", X"82", X"c0", X"07", X"c0", X"06", X"12", X"1a", 
    X"3e", X"d0", X"06", X"d0", X"07", X"80", X"db", X"90", 
    X"06", X"80", X"e0", X"ff", X"90", X"06", X"82", X"e0", 
    X"fd", X"c3", X"9f", X"50", X"09", X"90", X"06", X"80", 
    X"ef", X"c3", X"9d", X"f0", X"80", X"0c", X"90", X"06", 
    X"80", X"e4", X"f0", X"80", X"05", X"90", X"06", X"80", 
    X"ee", X"f0", X"90", X"06", X"8a", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"90", X"06", X"82", X"e0", X"fd", X"8d", 
    X"03", X"1d", X"eb", X"60", X"3e", X"b2", X"0e", X"20", 
    X"0e", X"14", X"0e", X"be", X"00", X"01", X"0f", X"8e", 
    X"82", X"8f", X"83", X"e0", X"c4", X"54", X"0f", X"fb", 
    X"90", X"06", X"6f", X"f0", X"80", X"0e", X"8e", X"82", 
    X"8f", X"83", X"e0", X"fb", X"53", X"03", X"0f", X"90", 
    X"06", X"6f", X"eb", X"f0", X"90", X"06", X"6f", X"e0", 
    X"f5", X"82", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"12", X"1a", X"7b", X"d0", X"05", X"d0", X"06", X"d0", 
    X"07", X"80", X"bc", X"20", X"06", X"03", X"02", X"1b", 
    X"46", X"90", X"06", X"80", X"e0", X"ff", X"8f", X"06", 
    X"1f", X"ee", X"70", X"03", X"02", X"1b", X"46", X"75", 
    X"82", X"20", X"c0", X"07", X"12", X"1a", X"3e", X"d0", 
    X"07", X"80", X"eb", X"8c", X"82", X"12", X"1a", X"3e", 
    X"02", X"1b", X"46", X"90", X"06", X"70", X"e0", X"fe", 
    X"a3", X"e0", X"8e", X"82", X"f5", X"83", X"22", X"aa", 
    X"82", X"ab", X"83", X"12", X"22", X"4f", X"60", X"03", 
    X"a3", X"80", X"f8", X"c3", X"e5", X"82", X"9a", X"f5", 
    X"82", X"e5", X"83", X"9b", X"f5", X"83", X"22", X"20", 
    X"f7", X"14", X"30", X"f6", X"14", X"88", X"83", X"a8", 
    X"82", X"20", X"f5", X"07", X"e6", X"a8", X"83", X"75", 
    X"83", X"00", X"22", X"e2", X"80", X"f7", X"e4", X"93", 
    X"22", X"e0", X"22", X"75", X"82", X"00", X"22", X"64", 
    X"68", X"72", X"79", X"2e", X"72", X"65", X"73", X"00", 
    X"61", X"2b", X"00", X"43", X"61", X"6e", X"20", X"6e", 
    X"6f", X"74", X"20", X"6f", X"70", X"65", X"6e", X"20", 
    X"64", X"68", X"72", X"79", X"2e", X"72", X"65", X"73", 
    X"0a", X"0a", X"00", X"44", X"48", X"52", X"59", X"53", 
    X"54", X"4f", X"4e", X"45", X"20", X"50", X"52", X"4f", 
    X"47", X"52", X"41", X"4d", X"2c", X"20", X"53", X"4f", 
    X"4d", X"45", X"20", X"53", X"54", X"52", X"49", X"4e", 
    X"47", X"00", X"44", X"48", X"52", X"59", X"53", X"54", 
    X"4f", X"4e", X"45", X"20", X"50", X"52", X"4f", X"47", 
    X"52", X"41", X"4d", X"2c", X"20", X"31", X"27", X"53", 
    X"54", X"20", X"53", X"54", X"52", X"49", X"4e", X"47", 
    X"00", X"0a", X"00", X"44", X"68", X"72", X"79", X"73", 
    X"74", X"6f", X"6e", X"65", X"20", X"42", X"65", X"6e", 
    X"63", X"68", X"6d", X"61", X"72", X"6b", X"2c", X"20", 
    X"56", X"65", X"72", X"73", X"69", X"6f", X"6e", X"20", 
    X"32", X"2e", X"31", X"20", X"28", X"4c", X"61", X"6e", 
    X"67", X"75", X"61", X"67", X"65", X"3a", X"20", X"43", 
    X"29", X"0a", X"00", X"45", X"78", X"65", X"63", X"75", 
    X"74", X"69", X"6f", X"6e", X"20", X"73", X"74", X"61", 
    X"72", X"74", X"73", X"2c", X"20", X"25", X"64", X"20", 
    X"72", X"75", X"6e", X"73", X"20", X"74", X"68", X"72", 
    X"6f", X"75", X"67", X"68", X"20", X"44", X"68", X"72", 
    X"79", X"73", X"74", X"6f", X"6e", X"65", X"0a", X"00", 
    X"44", X"48", X"52", X"59", X"53", X"54", X"4f", X"4e", 
    X"45", X"20", X"50", X"52", X"4f", X"47", X"52", X"41", 
    X"4d", X"2c", X"20", X"32", X"27", X"4e", X"44", X"20", 
    X"53", X"54", X"52", X"49", X"4e", X"47", X"00", X"44", 
    X"48", X"52", X"59", X"53", X"54", X"4f", X"4e", X"45", 
    X"20", X"50", X"52", X"4f", X"47", X"52", X"41", X"4d", 
    X"2c", X"20", X"33", X"27", X"52", X"44", X"20", X"53", 
    X"54", X"52", X"49", X"4e", X"47", X"00", X"45", X"78", 
    X"65", X"63", X"75", X"74", X"69", X"6f", X"6e", X"20", 
    X"65", X"6e", X"64", X"73", X"0a", X"00", X"46", X"69", 
    X"6e", X"61", X"6c", X"20", X"76", X"61", X"6c", X"75", 
    X"65", X"73", X"20", X"6f", X"66", X"20", X"74", X"68", 
    X"65", X"20", X"76", X"61", X"72", X"69", X"61", X"62", 
    X"6c", X"65", X"73", X"20", X"75", X"73", X"65", X"64", 
    X"20", X"69", X"6e", X"20", X"74", X"68", X"65", X"20", 
    X"62", X"65", X"6e", X"63", X"68", X"6d", X"61", X"72", 
    X"6b", X"3a", X"0a", X"00", X"49", X"6e", X"74", X"5f", 
    X"47", X"6c", X"6f", X"62", X"3a", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"25", X"64", X"0a", X"00", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"73", X"68", X"6f", 
    X"75", X"6c", X"64", X"20", X"62", X"65", X"3a", X"20", 
    X"20", X"20", X"25", X"64", X"0a", X"00", X"42", X"6f", 
    X"6f", X"6c", X"5f", X"47", X"6c", X"6f", X"62", X"3a", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"25", X"64", X"0a", X"00", X"43", 
    X"68", X"5f", X"31", X"5f", X"47", X"6c", X"6f", X"62", 
    X"3a", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"25", X"63", X"0a", X"00", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"73", X"68", X"6f", X"75", X"6c", X"64", X"20", X"62", 
    X"65", X"3a", X"20", X"20", X"20", X"25", X"63", X"0a", 
    X"00", X"43", X"68", X"5f", X"32", X"5f", X"47", X"6c", 
    X"6f", X"62", X"3a", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"25", X"63", 
    X"0a", X"00", X"41", X"72", X"72", X"5f", X"31", X"5f", 
    X"47", X"6c", X"6f", X"62", X"5b", X"38", X"5d", X"3a", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"25", 
    X"64", X"0a", X"00", X"41", X"72", X"72", X"5f", X"32", 
    X"5f", X"47", X"6c", X"6f", X"62", X"5b", X"38", X"5d", 
    X"5b", X"37", X"5d", X"3a", X"20", X"20", X"20", X"20", 
    X"25", X"64", X"0a", X"00", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"73", X"68", X"6f", X"75", 
    X"6c", X"64", X"20", X"62", X"65", X"3a", X"20", X"20", 
    X"20", X"4e", X"75", X"6d", X"62", X"65", X"72", X"5f", 
    X"4f", X"66", X"5f", X"52", X"75", X"6e", X"73", X"20", 
    X"2b", X"20", X"31", X"30", X"0a", X"00", X"50", X"74", 
    X"72", X"5f", X"47", X"6c", X"6f", X"62", X"2d", X"3e", 
    X"0a", X"00", X"20", X"20", X"50", X"74", X"72", X"5f", 
    X"43", X"6f", X"6d", X"70", X"3a", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"25", 
    X"64", X"0a", X"00", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"73", X"68", X"6f", X"75", X"6c", 
    X"64", X"20", X"62", X"65", X"3a", X"20", X"20", X"20", 
    X"28", X"69", X"6d", X"70", X"6c", X"65", X"6d", X"65", 
    X"6e", X"74", X"61", X"74", X"69", X"6f", X"6e", X"2d", 
    X"64", X"65", X"70", X"65", X"6e", X"64", X"65", X"6e", 
    X"74", X"29", X"0a", X"00", X"20", X"20", X"44", X"69", 
    X"73", X"63", X"72", X"3a", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"25", X"64", X"0a", X"00", X"20", X"20", X"45", 
    X"6e", X"75", X"6d", X"5f", X"43", X"6f", X"6d", X"70", 
    X"3a", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"25", X"64", X"0a", X"00", X"20", X"20", 
    X"49", X"6e", X"74", X"5f", X"43", X"6f", X"6d", X"70", 
    X"3a", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"25", X"64", X"0a", X"00", X"20", 
    X"20", X"53", X"74", X"72", X"5f", X"43", X"6f", X"6d", 
    X"70", X"3a", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"25", X"73", X"0a", X"00", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"73", X"68", X"6f", X"75", X"6c", X"64", X"20", X"62", 
    X"65", X"3a", X"20", X"20", X"20", X"44", X"48", X"52", 
    X"59", X"53", X"54", X"4f", X"4e", X"45", X"20", X"50", 
    X"52", X"4f", X"47", X"52", X"41", X"4d", X"2c", X"20", 
    X"53", X"4f", X"4d", X"45", X"20", X"53", X"54", X"52", 
    X"49", X"4e", X"47", X"0a", X"00", X"4e", X"65", X"78", 
    X"74", X"5f", X"50", X"74", X"72", X"5f", X"47", X"6c", 
    X"6f", X"62", X"2d", X"3e", X"0a", X"00", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"73", X"68", 
    X"6f", X"75", X"6c", X"64", X"20", X"62", X"65", X"3a", 
    X"20", X"20", X"20", X"28", X"69", X"6d", X"70", X"6c", 
    X"65", X"6d", X"65", X"6e", X"74", X"61", X"74", X"69", 
    X"6f", X"6e", X"2d", X"64", X"65", X"70", X"65", X"6e", 
    X"64", X"65", X"6e", X"74", X"29", X"2c", X"20", X"73", 
    X"61", X"6d", X"65", X"20", X"61", X"73", X"20", X"61", 
    X"62", X"6f", X"76", X"65", X"0a", X"00", X"49", X"6e", 
    X"74", X"5f", X"31", X"5f", X"4c", X"6f", X"63", X"3a", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"25", X"64", X"0a", X"00", X"49", 
    X"6e", X"74", X"5f", X"32", X"5f", X"4c", X"6f", X"63", 
    X"3a", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"25", X"64", X"0a", X"00", 
    X"49", X"6e", X"74", X"5f", X"33", X"5f", X"4c", X"6f", 
    X"63", X"3a", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"25", X"64", X"0a", 
    X"00", X"45", X"6e", X"75", X"6d", X"5f", X"4c", X"6f", 
    X"63", X"3a", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"25", X"64", 
    X"0a", X"00", X"53", X"74", X"72", X"5f", X"31", X"5f", 
    X"4c", X"6f", X"63", X"3a", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"25", 
    X"73", X"0a", X"00", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"73", X"68", X"6f", X"75", X"6c", 
    X"64", X"20", X"62", X"65", X"3a", X"20", X"20", X"20", 
    X"44", X"48", X"52", X"59", X"53", X"54", X"4f", X"4e", 
    X"45", X"20", X"50", X"52", X"4f", X"47", X"52", X"41", 
    X"4d", X"2c", X"20", X"31", X"27", X"53", X"54", X"20", 
    X"53", X"54", X"52", X"49", X"4e", X"47", X"0a", X"00", 
    X"53", X"74", X"72", X"5f", X"32", X"5f", X"4c", X"6f", 
    X"63", X"3a", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"25", X"73", X"0a", 
    X"00", X"20", X"20", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"73", X"68", X"6f", X"75", X"6c", X"64", X"20", 
    X"62", X"65", X"3a", X"20", X"20", X"20", X"44", X"48", 
    X"52", X"59", X"53", X"54", X"4f", X"4e", X"45", X"20", 
    X"50", X"52", X"4f", X"47", X"52", X"41", X"4d", X"2c", 
    X"20", X"32", X"27", X"4e", X"44", X"20", X"53", X"54", 
    X"52", X"49", X"4e", X"47", X"0a", X"00", X"54", X"69", 
    X"6d", X"65", X"20", X"65", X"6c", X"61", X"70", X"73", 
    X"65", X"64", X"3a", X"20", X"20", X"20", X"20", X"20", 
    X"20", X"20", X"20", X"20", X"20", X"25", X"6c", X"75", 
    X"2e", X"25", X"30", X"33", X"6c", X"75", X"20", X"73", 
    X"65", X"63", X"6f", X"6e", X"64", X"73", X"0a", X"00", 
    X"44", X"68", X"72", X"79", X"73", X"74", X"6f", X"6e", 
    X"65", X"73", X"20", X"70", X"65", X"72", X"20", X"73", 
    X"65", X"63", X"6f", X"6e", X"64", X"3a", X"20", X"25", 
    X"64", X"0a", X"0a", X"00", X"54", X"65", X"73", X"74", 
    X"20", X"66", X"69", X"6e", X"69", X"73", X"68", X"65", 
    X"64", X"2e", X"0a", X"0a", X"00", X"52", X"65", X"67", 
    X"69", X"73", X"74", X"65", X"72", X"20", X"6f", X"70", 
    X"74", X"69", X"6f", X"6e", X"20", X"73", X"65", X"6c", 
    X"65", X"63", X"74", X"65", X"64", X"2e", X"00", X"3c", 
    X"4e", X"4f", X"20", X"46", X"4c", X"4f", X"41", X"54", 
    X"3e", X"00", X"52", X"65", X"67", X"69", X"73", X"74", 
    X"65", X"72", X"20", X"6f", X"70", X"74", X"69", X"6f", 
    X"6e", X"20", X"73", X"65", X"6c", X"65", X"63", X"74", 
    X"65", X"64", X"2e", X"00" 
);


end package obj_code_pkg;
